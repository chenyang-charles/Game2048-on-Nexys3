`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    21:08:14 01/02/2015 
// Design Name: 
// Module Name:    move_event 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module move_event(
			input wire clk,
			input wire [15:0] xkey,
			input wire [4:0] btn,
			output reg win,
			output reg isEnd,
			output reg [63:0] map
    );

	parameter test_map = {
		16'b0000_0001_0010_0011,
		16'b0100_0101_0110_0111,
		16'b1000_1001_1010_1011,
		16'b0000_0000_0000_0000
	};
	
	parameter init_map = {
		16'b0001_0000_0000_0000,
		16'b0000_0000_0000_0000,
		16'b0000_0000_0000_0000,
		16'b0000_0000_0000_0000
	};

	reg clr, up, down, left, right;


	initial
	begin
		win <= 0;
		isEnd <= 0;
		map <= init_map;
		clr <= 0;
		up <= 0;
		down <= 0;
		left <= 0;
		right <= 0;
	end
		
	always @(posedge clk)
	begin
		if (xkey == 16'hf076 && btn[0] == 0)
		begin
			clr <= 0;
		end
		else if (xkey[7:0] == 8'h76 || btn[0] == 1)
		begin
			clr <= 1;
		end
		else
		begin
			clr <= 0;
		end
		
		if (xkey == 16'hf075 && btn[1] == 0)
		begin
			up <= 0;
		end
		else if (xkey[7:0] == 8'h75 || btn[1] == 1)
		begin
			up <= 1;
		end
		else
		begin
			up <= 0;
		end
		
		if (xkey == 16'hf06b && btn[2] == 0)
		begin
			left <= 0;
		end
		else if (xkey[7:0] == 8'h6b || btn[2] == 1)
		begin
			left <= 1;
		end
		else
		begin
			left <= 0;
		end
		
		if (xkey == 16'hf072 && btn[3] == 0)
		begin
			down <= 0;
		end
		else if (xkey[7:0] == 8'h72 || btn[3] == 1)
		begin
			down <= 1;
		end
		else
		begin
			down <= 0;
		end
		
		if (xkey == 16'hf074 && btn[4] == 0)
		begin
			right <= 0;
		end
		else if (xkey[7:0] == 8'h74 || btn[4] == 1)
		begin
			right <= 1;
		end
		else
		begin
			right <= 0;
		end
	end
	
	always @(posedge clk)
	begin
		if (clr == 1)
		begin
			win <= 0;
			isEnd <= 0;
			map <= init_map;
		end
		else
		if (up == 1)
		begin
			/*Up*/
			/*First line*/
			if (map[63:60] > 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0)
			begin
				map[15:12] <= map[63:60];
				map[63:60] <= 1;
			end
			else if (map[63:60] > 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
			begin
				if (map[15:12] == map[63:60])
				begin
					map[15:12] <= (map[63:60] + 1);
					map[63:60] <= 1;
				end
				else
				begin
					map[31:28] <= map[63:60];
					map[63:60] <= 1;
				end
			end
			else if (map[63:60] > 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] == 0)
			begin
				if (map[31:28] == map[63:60])
				begin
					map[15:12] <= (map[63:60] + 1);
					map[63:60] <= 0;
					map[31:28] <= 1;
				end
				else
				begin
					map[15:12] <= map[31:28];
					map[31:28] <= map[63:60];
					map[63:60] <= 1;
				end
			end
			else if (map[63:60] > 0 && map[47:44] > 0 && map[31:28] == 0 && map[15:12] == 0)
			begin
				if (map[47:44] == map[63:60])
				begin
					map[15:12] <= (map[63:60] + 1);
					map[63:60] <= 0;
					map[47:44] <= 1;
				end
				else
				begin
					map[15:12] <= map[47:44];
					map[31:28] <= map[63:60];
					map[47:44] <= 1;
					map[63:60] <= 0;
				end
			end
			else if (map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] == 0)
			begin
				if (map[31:28] == map[47:44])
				begin
					map[15:12] <= (map[31:28] + 1);
					map[31:28] <= map[63:60];
					map[63:60] <= 1;
					map[47:44] <= 0;
				end
				else
				if (map[63:60] == map[47:44])
				begin
					map[15:12] <= map[31:28];
					map[31:28] <= (map[47:44] + 1);
					map[63:60] <= 1;
					map[47:44] <= 0;
				end
				else
				begin
					map[15:12] <= map[31:28];
					map[31:28] <= map[47:44];
					map[63:60] <= 1;
					map[47:44] <= map[63:60];
				end
			end
			else if (map[63:60] > 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0)
			begin
				if (map[31:28] == map[15:12])
				begin
					map[15:12] <= (map[15:12] + 1);
					map[31:28] <= map[63:60];
					map[47:44] <= 1;
					map[63:60] <= 0;
				end
				else
				if (map[63:60] == map[31:28])
				begin
					map[31:28] <= (map[31:28] + 1);
					map[63:60] <= 1;
				end
				else
				begin
					map[47:44] <= map[63:60];
					map[63:60] <= 1;
				end
			end
			else if (map[63:60] > 0 && map[47:44] > 0 && map[31:28] == 0 && map[15:12] > 0)
			begin
				if (map[47:44] == map[15:12])
				begin
					map[15:12] <= (map[15:12] + 1);
					map[31:28] <= map[63:60];
					map[47:44] <= 0;
					map[63:60] <= 1;
				end
				else
				if (map[63:60] == map[47:44])
				begin
					map[31:28] <= (map[47:44] + 1);
					map[63:60] <= 1;
					map[47:44] <= 0;
				end
				else
				begin
					map[31:28] <= map[47:44];
					map[47:44] <= map[63:60];
					map[63:60] <= 1;
				end
			end
			else if (map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0)
			begin
				if (map[31:28] == map[15:12])
				begin
					map[15:12] <= (map[15:12] + 1);
					if (map[63:60] == map[47:44])
					begin
						map[31:28] <= (map[47:44] + 1);
						map[63:60] <= 1;
						map[47:44] <= 0;
					end
					else
					begin
						map[31:28] <= map[47:44];
						map[63:60] <= 1;
						map[47:44] <= map[63:60];
					end
				end
				else
				if (map[47:44] == map[31:28])
				begin
					map[31:28] <= (map[31:28] + 1);
					map[47:44] <= map[63:60];
					map[63:60] <= 1;
				end
				else
				if (map[63:60] == map[47:44])
				begin
					map[47:44] <= (map[47:44] + 1);
					map[63:60] <= 1;
				end
			end
			else if (map[63:60] == 0 && map[47:44] > 0 && map[31:28] == 0 && map[15:12] == 0)
			begin
				map[15:12] <= map[47:44];
				map[47:44] <= 1;
			end
			else if (map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] == 0)
			begin
				map[15:12] <= map[31:28];
				map[31:28] <= 1;
			end
			else if (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
			begin
			end
			else if (map[63:60] == 0 && map[47:44] > 0 && map[31:28] == 0 && map[15:12] > 0)
			begin
				if (map[15:12] == map[47:44])
				begin
					map[15:12] <= (map[15:12] + 1);
					map[47:44] <= 1;
				end
				else
				begin
					map[31:28] <= map[47:44];
					map[47:44] <= 1;
				end
			end
			else if (map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0)
			begin
				if (map[31:28] == map[15:12])
				begin
					map[15:12] <= (map[15:12] + 1);
					map[31:28] <= 1;
				end
			end
			else if (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] == 0)
			begin
				if (map[47:44] == map[31:28])
				begin
					map[15:12] <= (map[31:28] + 1);
					map[31:28] <= 0;
					map[47:44] <= 1;
				end
				else
				begin
					map[15:12] <= map[31:28];
					map[31:28] <= map[47:44];
					map[47:44] <= 1;
				end
			end
			else if (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0)
			begin
				if (map[15:12] == map[31:28])
				begin
					map[15:12] <= (map[31:28] + 1);
					map[31:28] <= map[47:44];
					map[47:44] <= 1;
				end
				else
				if (map[31:28] == map[47:44])
				begin
					map[31:28] <= (map[31:28] + 1);
					map[47:44] <= 1;
				end
			end
			else if (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0)
			begin
			end
			
			/*Second line*/			
			
			if (map[59:56] > 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0)
			begin
				map[11:8] <= map[59:56];
				if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
				begin
					map[59:56] <= 1;
				end
				else
				begin
					map[59:56] <= 0;
				end
			end
			else if (map[59:56] > 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
			begin
				if (map[11:8] == map[59:56])
				begin
					map[11:8] <= (map[59:56] + 1);
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
				else
				begin
					map[27:24] <= map[59:56];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
			end
			else if (map[59:56] > 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] == 0)
			begin
				if (map[27:24] == map[59:56])
				begin
					map[11:8] <= (map[59:56] + 1);
					map[59:56] <= 0;
					map[27:24] <= 1;
				end
				else
				begin
					map[11:8] <= map[27:24];
					map[27:24] <= map[59:56];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
			end
			else if (map[59:56] > 0 && map[43:40] > 0 && map[27:24] == 0 && map[11:8] == 0)
			begin
				if (map[43:40] == map[59:56])
				begin
					map[11:8] <= (map[59:56] + 1);
					map[59:56] <= 0;
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
					   	map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
				else
				begin
					map[11:8] <= map[43:40];
					map[27:24] <= map[59:56];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
					map[59:56] <= 0;
				end
			end
			else if (map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] == 0)
			begin
				if (map[27:24] == map[43:40])
				begin
					map[11:8] <= (map[27:24] + 1);
					map[27:24] <= map[59:56];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
					map[43:40] <= 0;
				end
				else
				if (map[59:56] == map[43:40])
				begin
					map[11:8] <= map[27:24];
					map[27:24] <= (map[43:40] + 1);
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
					map[43:40] <= 0;
				end
				else
				begin
					map[11:8] <= map[27:24];
					map[27:24] <= map[43:40];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
					map[43:40] <= map[59:56];
				end
			end
			else if (map[59:56] > 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0)
			begin
				if (map[27:24] == map[11:8])
				begin
					map[11:8] <= (map[11:8] + 1);
					map[27:24] <= map[59:56];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
					    map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
					map[59:56] <= 0;
				end
				else
				if (map[59:56] == map[27:24])
				begin
					map[27:24] <= (map[27:24] + 1);
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
				else
				begin
					map[43:40] <= map[59:56];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
			end
			else if (map[59:56] > 0 && map[43:40] > 0 && map[27:24] == 0 && map[11:8] > 0)
			begin
				if (map[43:40] == map[11:8])
				begin
					map[11:8] <= (map[11:8] + 1);
					map[27:24] <= map[59:56];
					map[43:40] <= 0;
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
				else
				if (map[59:56] == map[43:40])
				begin
					map[27:24] <= (map[43:40] + 1);
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
					map[43:40] <= 0;
				end
				else
				begin
					map[27:24] <= map[43:40];
					map[43:40] <= map[59:56];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
			end
			else if (map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0)
			begin
				if (map[27:24] == map[11:8])
				begin
					map[11:8] <= (map[11:8] + 1);
					if (map[59:56] == map[43:40])
					begin
						map[27:24] <= (map[43:40] + 1);
						if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
						begin
							map[59:56] <= 1;
						end
						else
						begin
							map[59:56] <= 0;
						end
						map[43:40] <= 0;
					end
					else
					begin
						map[27:24] <= map[43:40];
						if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
						begin
							map[59:56] <= 1;
						end
						else
						begin
							map[59:56] <= 0;
						end
						map[43:40] <= map[59:56];
					end
				end
				else
				if (map[43:40] == map[27:24])
				begin
					map[27:24] <= (map[27:24] + 1);
					map[43:40] <= map[59:56];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
				else
				if (map[59:56] == map[43:40])
				begin
					map[43:40] <= (map[43:40] + 1);
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
			end
			else if (map[59:56] == 0 && map[43:40] > 0 && map[27:24] == 0 && map[11:8] == 0)
			begin
				map[11:8] <= map[43:40];
				if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
				begin
					map[43:40] <= 1;
				end
				else
				begin
					map[43:40] <= 0;
				end
			end
			else if (map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] == 0)
			begin
				map[11:8] <= map[27:24];
				map[27:24] <= 1;
			end
			else if (map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
			begin
			end
			else if (map[59:56] == 0 && map[43:40] > 0 && map[27:24] == 0 && map[11:8] > 0)
			begin
				if (map[11:8] == map[43:40])
				begin
					map[11:8] <= (map[11:8] + 1);
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
				else
				begin
					map[27:24] <= map[43:40];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
			end
			else if (map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0)
			begin
				if (map[27:24] == map[11:8])
				begin
					map[11:8] <= (map[11:8] + 1);
					map[27:24] <= 1;
				end
			end
			else if (map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] == 0)
			begin
				if (map[43:40] == map[27:24])
				begin
					map[11:8] <= (map[27:24] + 1);
					map[27:24] <= 0;
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
				else
				begin
					map[11:8] <= map[27:24];
					map[27:24] <= map[43:40];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
			end
			else if (map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0)
			begin
				if (map[11:8] == map[27:24])
				begin
					map[11:8] <= (map[27:24] + 1);
					map[27:24] <= map[43:40];
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
				else
				if (map[27:24] == map[43:40])
				begin
					map[27:24] <= (map[27:24] + 1);
					if ((map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0
				&& map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || (map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
				(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || (map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0))
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
			end
			else if (map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0)
			begin
			end

			/*Third line*/			
			
			if (map[55:52] > 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0)
			begin
				map[7:4] <= map[55:52];
				if 
				( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
				begin
					map[55:52] <= 1;
				end
				else
				begin
					map[55:52] <= 0;
				end
			end
			else if (map[55:52] > 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
			begin
				if (map[7:4] == map[55:52])
				begin
					map[7:4] <= (map[55:52] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
				else
				begin
					map[23:20] <= map[55:52];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
			end
			else if (map[55:52] > 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] == 0)
			begin
				if (map[23:20] == map[55:52])
				begin
					map[7:4] <= (map[55:52] + 1);
					map[55:52] <= 0;
					map[23:20] <= 1;
				end
				else
				begin
					map[7:4] <= map[23:20];
					map[23:20] <= map[55:52];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
			end
			else if (map[55:52] > 0 && map[39:36] > 0 && map[23:20] == 0 && map[7:4] == 0)
			begin
				if (map[39:36] == map[55:52])
				begin
					map[7:4] <= (map[55:52] + 1);
					map[55:52] <= 0;
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
					   	map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
				else
				begin
					map[7:4] <= map[39:36];
					map[23:20] <= map[55:52];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
					map[55:52] <= 0;
				end
			end
			else if (map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] == 0)
			begin
				if (map[23:20] == map[39:36])
				begin
					map[7:4] <= (map[23:20] + 1);
					map[23:20] <= map[55:52];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
					map[39:36] <= 0;
				end
				else
				if (map[55:52] == map[39:36])
				begin
					map[7:4] <= map[23:20];
					map[23:20] <= (map[39:36] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
					map[39:36] <= 0;
				end
				else
				begin
					map[7:4] <= map[23:20];
					map[23:20] <= map[39:36];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
					map[39:36] <= map[55:52];
				end
			end
			else if (map[55:52] > 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0)
			begin
				if (map[23:20] == map[7:4])
				begin
					map[7:4] <= (map[7:4] + 1);
					map[23:20] <= map[55:52];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
					    map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
					map[55:52] <= 0;
				end
				else
				if (map[55:52] == map[23:20])
				begin
					map[23:20] <= (map[23:20] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
				else
				begin
					map[39:36] <= map[55:52];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
			end
			else if (map[55:52] > 0 && map[39:36] > 0 && map[23:20] == 0 && map[7:4] > 0)
			begin
				if (map[39:36] == map[7:4])
				begin
					map[7:4] <= (map[7:4] + 1);
					map[23:20] <= map[55:52];
					map[39:36] <= 0;
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
				else
				if (map[55:52] == map[39:36])
				begin
					map[23:20] <= (map[39:36] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
					map[39:36] <= 0;
				end
				else
				begin
					map[23:20] <= map[39:36];
					map[39:36] <= map[55:52];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
			end
			else if (map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0)
			begin
				if (map[23:20] == map[7:4])
				begin
					map[7:4] <= (map[7:4] + 1);
					if (map[55:52] == map[39:36])
					begin
						map[23:20] <= (map[39:36] + 1);
						if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
						begin
							map[55:52] <= 1;
						end
						else
						begin
							map[55:52] <= 0;
						end
						map[39:36] <= 0;
					end
					else
					begin
						map[23:20] <= map[39:36];
						if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
						begin
							map[55:52] <= 1;
						end
						else
						begin
							map[55:52] <= 0;
						end
						map[39:36] <= map[55:52];
					end
				end
				else
				if (map[39:36] == map[23:20])
				begin
					map[23:20] <= (map[23:20] + 1);
					map[39:36] <= map[55:52];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
				else
				if (map[55:52] == map[39:36])
				begin
					map[39:36] <= (map[39:36] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
			end
			else if (map[55:52] == 0 && map[39:36] > 0 && map[23:20] == 0 && map[7:4] == 0)
			begin
				map[7:4] <= map[39:36];
				if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
				begin
					map[39:36] <= 1;
				end
				else
				begin
					map[39:36] <= 0;
				end
			end
			else if (map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] == 0)
			begin
				map[7:4] <= map[23:20];
				map[23:20] <= 1;
			end
			else if (map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
			begin
			end
			else if (map[55:52] == 0 && map[39:36] > 0 && map[23:20] == 0 && map[7:4] > 0)
			begin
				if (map[7:4] == map[39:36])
				begin
					map[7:4] <= (map[7:4] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
				else
				begin
					map[23:20] <= map[39:36];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
			end
			else if (map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0)
			begin
				if (map[23:20] == map[7:4])
				begin
					map[7:4] <= (map[7:4] + 1);
					map[23:20] <= 1;
				end
			end
			else if (map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] == 0)
			begin
				if (map[39:36] == map[23:20])
				begin
					map[7:4] <= (map[23:20] + 1);
					map[23:20] <= 0;
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
				else
				begin
					map[7:4] <= map[23:20];
					map[23:20] <= map[39:36];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
			end
			else if (map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0)
			begin
				if (map[7:4] == map[23:20])
				begin
					map[7:4] <= (map[23:20] + 1);
					map[23:20] <= map[39:36];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
				else
				if (map[23:20] == map[39:36])
				begin
					map[23:20] <= (map[23:20] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
			end
			else if (map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0)
			begin
			end

			/*Forth line*/			
			
			if (map[51:48] > 0 && map[35:32] == 0 && map[19:16] == 0 && map[3:0] == 0)
			begin
				map[3:0] <= map[51:48];
				if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
				begin
					map[51:48] <= 1;
				end
				else
				begin
					map[51:48] <= 0;
				end
			end
			else if (map[51:48] > 0 && map[35:32] == 0 && map[19:16] == 0 && map[3:0] > 0)
			begin
				if (map[3:0] == map[51:48])
				begin
					map[3:0] <= (map[51:48] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
				else
				begin
					map[19:16] <= map[51:48];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] > 0 && map[35:32] == 0 && map[19:16] > 0 && map[3:0] == 0)
			begin
				if (map[19:16] == map[51:48])
				begin
					map[3:0] <= (map[51:48] + 1);
					map[51:48] <= 0;
					map[19:16] <= 1;
				end
				else
				begin
					map[3:0] <= map[19:16];
					map[19:16] <= map[51:48];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] > 0 && map[35:32] > 0 && map[19:16] == 0 && map[3:0] == 0)
			begin
				if (map[35:32] == map[51:48])
				begin
					map[3:0] <= (map[51:48] + 1);
					map[51:48] <= 0;
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
					   	map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
				else
				begin
					map[3:0] <= map[35:32];
					map[19:16] <= map[51:48];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
					map[51:48] <= 0;
				end
			end
			else if (map[51:48] > 0 && map[35:32] > 0 && map[19:16] > 0 && map[3:0] == 0)
			begin
				if (map[19:16] == map[35:32])
				begin
					map[3:0] <= (map[19:16] + 1);
					map[19:16] <= map[51:48];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
					map[35:32] <= 0;
				end
				else
				if (map[51:48] == map[35:32])
				begin
					map[3:0] <= map[19:16];
					map[19:16] <= (map[35:32] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
					map[35:32] <= 0;
				end
				else
				begin
					map[3:0] <= map[19:16];
					map[19:16] <= map[35:32];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
					map[35:32] <= map[51:48];
				end
			end
			else if (map[51:48] > 0 && map[35:32] == 0 && map[19:16] > 0 && map[3:0] > 0)
			begin
				if (map[19:16] == map[3:0])
				begin
					map[3:0] <= (map[3:0] + 1);
					map[19:16] <= map[51:48];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
					    map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
					map[51:48] <= 0;
				end
				else
				if (map[51:48] == map[19:16])
				begin
					map[19:16] <= (map[19:16] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
				else
				begin
					map[35:32] <= map[51:48];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] > 0 && map[35:32] > 0 && map[19:16] == 0 && map[3:0] > 0)
			begin
				if (map[35:32] == map[3:0])
				begin
					map[3:0] <= (map[3:0] + 1);
					map[19:16] <= map[51:48];
					map[35:32] <= 0;
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
				else
				if (map[51:48] == map[35:32])
				begin
					map[19:16] <= (map[35:32] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
					map[35:32] <= 0;
				end
				else
				begin
					map[19:16] <= map[35:32];
					map[35:32] <= map[51:48];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] > 0 && map[35:32] > 0 && map[19:16] > 0 && map[3:0] > 0)
			begin
				if (map[19:16] == map[3:0])
				begin
					map[3:0] <= (map[3:0] + 1);
					if (map[51:48] == map[35:32])
					begin
						map[19:16] <= (map[35:32] + 1);
						if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
						begin
							map[51:48] <= 1;
						end
						else
						begin
							map[51:48] <= 0;
						end
						map[35:32] <= 0;
					end
					else
					begin
						map[19:16] <= map[35:32];
						if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
						begin
							map[51:48] <= 1;
						end
						else
						begin
							map[51:48] <= 0;
						end
						map[35:32] <= map[51:48];
					end
				end
				else
				if (map[35:32] == map[19:16])
				begin
					map[19:16] <= (map[19:16] + 1);
					map[35:32] <= map[51:48];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
				else
				if (map[51:48] == map[35:32])
				begin
					map[35:32] <= (map[35:32] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] == 0 && map[35:32] > 0 && map[19:16] == 0 && map[3:0] == 0)
			begin
				map[3:0] <= map[35:32];
				if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
				begin
					map[35:32] <= 1;
				end
				else
				begin
					map[35:32] <= 0;
				end
			end
			else if (map[51:48] == 0 && map[35:32] == 0 && map[19:16] > 0 && map[3:0] == 0)
			begin
				map[3:0] <= map[19:16];
				map[19:16] <= 1;
			end
			else if (map[51:48] == 0 && map[35:32] == 0 && map[19:16] == 0 && map[3:0] > 0)
			begin
			end
			else if (map[51:48] == 0 && map[35:32] > 0 && map[19:16] == 0 && map[3:0] > 0)
			begin
				if (map[3:0] == map[35:32])
				begin
					map[3:0] <= (map[3:0] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
				else
				begin
					map[19:16] <= map[35:32];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
			end
			else if (map[51:48] == 0 && map[35:32] == 0 && map[19:16] > 0 && map[3:0] > 0)
			begin
				if (map[19:16] == map[3:0])
				begin
					map[3:0] <= (map[3:0] + 1);
					map[19:16] <= 1;
				end
			end
			else if (map[51:48] == 0 && map[35:32] > 0 && map[19:16] > 0 && map[3:0] == 0)
			begin
				if (map[35:32] == map[19:16])
				begin
					map[3:0] <= (map[19:16] + 1);
					map[19:16] <= 0;
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
				else
				begin
					map[3:0] <= map[19:16];
					map[19:16] <= map[35:32];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
			end
			else if (map[51:48] == 0 && map[35:32] > 0 && map[19:16] > 0 && map[3:0] > 0)
			begin
				if (map[3:0] == map[19:16])
				begin
					map[3:0] <= (map[19:16] + 1);
					map[19:16] <= map[35:32];
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
				else
				if (map[19:16] == map[35:32])
				begin
					map[19:16] <= (map[19:16] + 1);
					if ( 
					( 
						(map[63:60] > 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[63:60] != map[47:44] && map[47:44] != map[31:28] && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] == 0) || 
						(map[63:60] == 0 && map[47:44] > 0 && map[31:28] > 0 && map[15:12] > 0 && map[47:44] != map[31:28] && map[31:28] != map[15:12]) ||
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] > 0 && map[15:12] > 0 && map[31:28] != map[15:12]) || 
						(map[63:60] == 0 && map[47:44] == 0 && map[31:28] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[59:56] > 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[59:56] != map[43:40] && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] == 0) || 
						(map[59:56] == 0 && map[43:40] > 0 && map[27:24] > 0 && map[11:8] > 0 && map[43:40] != map[27:24] && map[27:24] != map[11:8]) ||
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] > 0 && map[11:8] > 0 && map[27:24] != map[11:8]) || 
						(map[59:56] == 0 && map[43:40] == 0 && map[27:24] == 0 && map[11:8] > 0)
					)
					&& 
					(	
						(map[55:52] > 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[55:52] != map[39:36] && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] == 0) || 
						(map[55:52] == 0 && map[39:36] > 0 && map[23:20] > 0 && map[7:4] > 0 && map[39:36] != map[23:20] && map[23:20] != map[7:4]) ||
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] > 0 && map[7:4] > 0 && map[23:20] != map[7:4]) || 
						(map[55:52] == 0 && map[39:36] == 0 && map[23:20] == 0 && map[7:4] > 0)
					)
				)
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
			end
			else if (map[51:48] == 0 && map[35:32] == 0 && map[19:16] == 0 && map[3:0] == 0)
			begin
			end
		end
		else
		if (left == 1)
		begin
			/*Left*/
			/*First line*/
			if (map[15:12] > 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0)
			begin
				map[3:0] <= map[15:12];
				map[15:12] <= 1;
			end
			else if (map[15:12] > 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
			begin
				if (map[3:0] == map[15:12])
				begin
					map[3:0] <= (map[15:12] + 1);
					map[15:12] <= 1;
				end
				else
				begin
					map[7:4] <= map[15:12];
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] > 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] == 0)
			begin
				if (map[7:4] == map[15:12])
				begin
					map[3:0] <= (map[15:12] + 1);
					map[15:12] <= 0;
					map[7:4] <= 1;
				end
				else
				begin
					map[3:0] <= map[7:4];
					map[7:4] <= map[15:12];
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] > 0 && map[11:8] > 0 && map[7:4] == 0 && map[3:0] == 0)
			begin
				if (map[11:8] == map[15:12])
				begin
					map[3:0] <= (map[15:12] + 1);
					map[15:12] <= 0;
					map[11:8] <= 1;
				end
				else
				begin
					map[3:0] <= map[11:8];
					map[7:4] <= map[15:12];
					map[11:8] <= 1;
					map[15:12] <= 0;
				end
			end
			else if (map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] == 0)
			begin
				if (map[7:4] == map[11:8])
				begin
					map[3:0] <= (map[7:4] + 1);
					map[7:4] <= map[15:12];
					map[15:12] <= 1;
					map[11:8] <= 0;
				end
				else
				if (map[15:12] == map[11:8])
				begin
					map[3:0] <= map[7:4];
					map[7:4] <= (map[11:8] + 1);
					map[15:12] <= 1;
					map[11:8] <= 0;
				end
				else
				begin
					map[3:0] <= map[7:4];
					map[7:4] <= map[11:8];
					map[15:12] <= 1;
					map[11:8] <= map[15:12];
				end
			end
			else if (map[15:12] > 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0)
			begin
				if (map[7:4] == map[3:0])
				begin
					map[3:0] <= (map[3:0] + 1);
					map[7:4] <= map[15:12];
					map[11:8] <= 1;
					map[15:12] <= 0;
				end
				else
				if (map[15:12] == map[7:4])
				begin
					map[7:4] <= (map[7:4] + 1);
					map[15:12] <= 1;
				end
				else
				begin
					map[11:8] <= map[15:12];
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] > 0 && map[11:8] > 0 && map[7:4] == 0 && map[3:0] > 0)
			begin
				if (map[11:8] == map[3:0])
				begin
					map[3:0] <= (map[3:0] + 1);
					map[7:4] <= map[15:12];
					map[11:8] <= 0;
					map[15:12] <= 1;
				end
				else
				if (map[15:12] == map[11:8])
				begin
					map[7:4] <= (map[11:8] + 1);
					map[15:12] <= 1;
					map[11:8] <= 0;
				end
				else
				begin
					map[7:4] <= map[11:8];
					map[11:8] <= map[15:12];
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0)
			begin
				if (map[7:4] == map[3:0])
				begin
					map[3:0] <= (map[3:0] + 1);
					if (map[15:12] == map[11:8])
					begin
						map[7:4] <= (map[11:8] + 1);
						map[15:12] <= 1;
						map[11:8] <= 0;
					end
					else
					begin
						map[7:4] <= map[11:8];
						map[15:12] <= 1;
						map[11:8] <= map[15:12];
					end
				end
				else
				if (map[11:8] == map[7:4])
				begin
					map[7:4] <= (map[7:4] + 1);
					map[11:8] <= map[15:12];
					map[15:12] <= 1;
				end
				else
				if (map[15:12] == map[11:8])
				begin
					map[11:8] <= (map[11:8] + 1);
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[11:8] > 0 && map[7:4] == 0 && map[3:0] == 0)
			begin
				map[3:0] <= map[11:8];
				map[11:8] <= 1;
			end
			else if (map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] == 0)
			begin
				map[3:0] <= map[7:4];
				map[7:4] <= 1;
			end
			else if (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
			begin
			end
			else if (map[15:12] == 0 && map[11:8] > 0 && map[7:4] == 0 && map[3:0] > 0)
			begin
				if (map[3:0] == map[11:8])
				begin
					map[3:0] <= (map[3:0] + 1);
					map[11:8] <= 1;
				end
				else
				begin
					map[7:4] <= map[11:8];
					map[11:8] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0)
			begin
				if (map[7:4] == map[3:0])
				begin
					map[3:0] <= (map[3:0] + 1);
					map[7:4] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] == 0)
			begin
				if (map[11:8] == map[7:4])
				begin
					map[3:0] <= (map[7:4] + 1);
					map[7:4] <= 0;
					map[11:8] <= 1;
				end
				else
				begin
					map[3:0] <= map[7:4];
					map[7:4] <= map[11:8];
					map[11:8] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0)
			begin
				if (map[3:0] == map[7:4])
				begin
					map[3:0] <= (map[7:4] + 1);
					map[7:4] <= map[11:8];
					map[11:8] <= 1;
				end
				else
				if (map[7:4] == map[11:8])
				begin
					map[7:4] <= (map[7:4] + 1);
					map[11:8] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0)
			begin
			end
			
			/*Second line*/			
			
			if (map[31:28] > 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0)
			begin
				map[19:16] <= map[31:28];
				if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
				begin
					map[31:28] <= 1;
				end
				else
				begin
					map[31:28] <= 0;
				end
			end
			else if (map[31:28] > 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
			begin
				if (map[19:16] == map[31:28])
				begin
					map[19:16] <= (map[31:28] + 1);
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
				else
				begin
					map[23:20] <= map[31:28];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
			end
			else if (map[31:28] > 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] == 0)
			begin
				if (map[23:20] == map[31:28])
				begin
					map[19:16] <= (map[31:28] + 1);
					map[31:28] <= 0;
					map[23:20] <= 1;
				end
				else
				begin
					map[19:16] <= map[23:20];
					map[23:20] <= map[31:28];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
			end
			else if (map[31:28] > 0 && map[27:24] > 0 && map[23:20] == 0 && map[19:16] == 0)
			begin
				if (map[27:24] == map[31:28])
				begin
					map[19:16] <= (map[31:28] + 1);
					map[31:28] <= 0;
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
					   	map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
				else
				begin
					map[19:16] <= map[27:24];
					map[23:20] <= map[31:28];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
					map[31:28] <= 0;
				end
			end
			else if (map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] == 0)
			begin
				if (map[23:20] == map[27:24])
				begin
					map[19:16] <= (map[23:20] + 1);
					map[23:20] <= map[31:28];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
					map[27:24] <= 0;
				end
				else
				if (map[31:28] == map[27:24])
				begin
					map[19:16] <= map[23:20];
					map[23:20] <= (map[27:24] + 1);
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
					map[27:24] <= 0;
				end
				else
				begin
					map[19:16] <= map[23:20];
					map[23:20] <= map[27:24];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
					map[27:24] <= map[31:28];
				end
			end
			else if (map[31:28] > 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0)
			begin
				if (map[23:20] == map[19:16])
				begin
					map[19:16] <= (map[19:16] + 1);
					map[23:20] <= map[31:28];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
					    map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
					map[31:28] <= 0;
				end
				else
				if (map[31:28] == map[23:20])
				begin
					map[23:20] <= (map[23:20] + 1);
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
				else
				begin
					map[27:24] <= map[31:28];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
			end
			else if (map[31:28] > 0 && map[27:24] > 0 && map[23:20] == 0 && map[19:16] > 0)
			begin
				if (map[27:24] == map[19:16])
				begin
					map[19:16] <= (map[19:16] + 1);
					map[23:20] <= map[31:28];
					map[27:24] <= 0;
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
				else
				if (map[31:28] == map[27:24])
				begin
					map[23:20] <= (map[27:24] + 1);
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
					map[27:24] <= 0;
				end
				else
				begin
					map[23:20] <= map[27:24];
					map[27:24] <= map[31:28];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
			end
			else if (map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0)
			begin
				if (map[23:20] == map[19:16])
				begin
					map[19:16] <= (map[19:16] + 1);
					if (map[31:28] == map[27:24])
					begin
						map[23:20] <= (map[27:24] + 1);
						if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
						begin
							map[31:28] <= 1;
						end
						else
						begin
							map[31:28] <= 0;
						end
						map[27:24] <= 0;
					end
					else
					begin
						map[23:20] <= map[27:24];
						if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
						begin
							map[31:28] <= 1;
						end
						else
						begin
							map[31:28] <= 0;
						end
						map[27:24] <= map[31:28];
					end
				end
				else
				if (map[27:24] == map[23:20])
				begin
					map[23:20] <= (map[23:20] + 1);
					map[27:24] <= map[31:28];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
				else
				if (map[31:28] == map[27:24])
				begin
					map[27:24] <= (map[27:24] + 1);
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[31:28] <= 1;
					end
					else
					begin
						map[31:28] <= 0;
					end
				end
			end
			else if (map[31:28] == 0 && map[27:24] > 0 && map[23:20] == 0 && map[19:16] == 0)
			begin
				map[19:16] <= map[27:24];
				if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
				begin
					map[27:24] <= 1;
				end
				else
				begin
					map[27:24] <= 0;
				end
			end
			else if (map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] == 0)
			begin
				map[19:16] <= map[23:20];
				map[23:20] <= 1;
			end
			else if (map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
			begin
			end
			else if (map[31:28] == 0 && map[27:24] > 0 && map[23:20] == 0 && map[19:16] > 0)
			begin
				if (map[19:16] == map[27:24])
				begin
					map[19:16] <= (map[19:16] + 1);
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
				else
				begin
					map[23:20] <= map[27:24];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
			end
			else if (map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0)
			begin
				if (map[23:20] == map[19:16])
				begin
					map[19:16] <= (map[19:16] + 1);
					map[23:20] <= 1;
				end
			end
			else if (map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] == 0)
			begin
				if (map[27:24] == map[23:20])
				begin
					map[19:16] <= (map[23:20] + 1);
					map[23:20] <= 0;
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
				else
				begin
					map[19:16] <= map[23:20];
					map[23:20] <= map[27:24];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
			end
			else if (map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0)
			begin
				if (map[19:16] == map[23:20])
				begin
					map[19:16] <= (map[23:20] + 1);
					map[23:20] <= map[27:24];
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
				else
				if (map[23:20] == map[27:24])
				begin
					map[23:20] <= (map[23:20] + 1);
					if ((map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0
				&& map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || (map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
				(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || (map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
			end
			else if (map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0)
			begin
			end

			/*Third line*/			
			
			if (map[47:44] > 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0)
			begin
				map[35:32] <= map[47:44];
				if 
				( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
				begin
					map[47:44] <= 1;
				end
				else
				begin
					map[47:44] <= 0;
				end
			end
			else if (map[47:44] > 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
			begin
				if (map[35:32] == map[47:44])
				begin
					map[35:32] <= (map[47:44] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
				else
				begin
					map[39:36] <= map[47:44];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
			end
			else if (map[47:44] > 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] == 0)
			begin
				if (map[39:36] == map[47:44])
				begin
					map[35:32] <= (map[47:44] + 1);
					map[47:44] <= 0;
					map[39:36] <= 1;
				end
				else
				begin
					map[35:32] <= map[39:36];
					map[39:36] <= map[47:44];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
			end
			else if (map[47:44] > 0 && map[43:40] > 0 && map[39:36] == 0 && map[35:32] == 0)
			begin
				if (map[43:40] == map[47:44])
				begin
					map[35:32] <= (map[47:44] + 1);
					map[47:44] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
					   	map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
				else
				begin
					map[35:32] <= map[43:40];
					map[39:36] <= map[47:44];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
					map[47:44] <= 0;
				end
			end
			else if (map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] == 0)
			begin
				if (map[39:36] == map[43:40])
				begin
					map[35:32] <= (map[39:36] + 1);
					map[39:36] <= map[47:44];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
					map[43:40] <= 0;
				end
				else
				if (map[47:44] == map[43:40])
				begin
					map[35:32] <= map[39:36];
					map[39:36] <= (map[43:40] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
					map[43:40] <= 0;
				end
				else
				begin
					map[35:32] <= map[39:36];
					map[39:36] <= map[43:40];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
					map[43:40] <= map[47:44];
				end
			end
			else if (map[47:44] > 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0)
			begin
				if (map[39:36] == map[35:32])
				begin
					map[35:32] <= (map[35:32] + 1);
					map[39:36] <= map[47:44];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
					    map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
					map[47:44] <= 0;
				end
				else
				if (map[47:44] == map[39:36])
				begin
					map[39:36] <= (map[39:36] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
				else
				begin
					map[43:40] <= map[47:44];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
			end
			else if (map[47:44] > 0 && map[43:40] > 0 && map[39:36] == 0 && map[35:32] > 0)
			begin
				if (map[43:40] == map[35:32])
				begin
					map[35:32] <= (map[35:32] + 1);
					map[39:36] <= map[47:44];
					map[43:40] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
				else
				if (map[47:44] == map[43:40])
				begin
					map[39:36] <= (map[43:40] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
					map[43:40] <= 0;
				end
				else
				begin
					map[39:36] <= map[43:40];
					map[43:40] <= map[47:44];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
			end
			else if (map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0)
			begin
				if (map[39:36] == map[35:32])
				begin
					map[35:32] <= (map[35:32] + 1);
					if (map[47:44] == map[43:40])
					begin
						map[39:36] <= (map[43:40] + 1);
						if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
						begin
							map[47:44] <= 1;
						end
						else
						begin
							map[47:44] <= 0;
						end
						map[43:40] <= 0;
					end
					else
					begin
						map[39:36] <= map[43:40];
						if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
						begin
							map[47:44] <= 1;
						end
						else
						begin
							map[47:44] <= 0;
						end
						map[43:40] <= map[47:44];
					end
				end
				else
				if (map[43:40] == map[39:36])
				begin
					map[39:36] <= (map[39:36] + 1);
					map[43:40] <= map[47:44];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
				else
				if (map[47:44] == map[43:40])
				begin
					map[43:40] <= (map[43:40] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[47:44] <= 1;
					end
					else
					begin
						map[47:44] <= 0;
					end
				end
			end
			else if (map[47:44] == 0 && map[43:40] > 0 && map[39:36] == 0 && map[35:32] == 0)
			begin
				map[35:32] <= map[43:40];
				if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
				begin
					map[43:40] <= 1;
				end
				else
				begin
					map[43:40] <= 0;
				end
			end
			else if (map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] == 0)
			begin
				map[35:32] <= map[39:36];
				map[39:36] <= 1;
			end
			else if (map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
			begin
			end
			else if (map[47:44] == 0 && map[43:40] > 0 && map[39:36] == 0 && map[35:32] > 0)
			begin
				if (map[35:32] == map[43:40])
				begin
					map[35:32] <= (map[35:32] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
				else
				begin
					map[39:36] <= map[43:40];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
			end
			else if (map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0)
			begin
				if (map[39:36] == map[35:32])
				begin
					map[35:32] <= (map[35:32] + 1);
					map[39:36] <= 1;
				end
			end
			else if (map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] == 0)
			begin
				if (map[43:40] == map[39:36])
				begin
					map[35:32] <= (map[39:36] + 1);
					map[39:36] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
				else
				begin
					map[35:32] <= map[39:36];
					map[39:36] <= map[43:40];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
			end
			else if (map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0)
			begin
				if (map[35:32] == map[39:36])
				begin
					map[35:32] <= (map[39:36] + 1);
					map[39:36] <= map[43:40];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
				else
				if (map[39:36] == map[43:40])
				begin
					map[39:36] <= (map[39:36] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
				)	
					begin
						map[43:40] <= 1;
					end
					else
					begin
						map[43:40] <= 0;
					end
				end
			end
			else if (map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0)
			begin
			end

			/*Forth line*/			
			
			if (map[63:60] > 0 && map[59:56] == 0 && map[55:52] == 0 && map[51:48] == 0)
			begin
				map[51:48] <= map[63:60];
				if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
				begin
					map[63:60] <= 1;
				end
				else
				begin
					map[63:60] <= 0;
				end
			end
			else if (map[63:60] > 0 && map[59:56] == 0 && map[55:52] == 0 && map[51:48] > 0)
			begin
				if (map[51:48] == map[63:60])
				begin
					map[51:48] <= (map[63:60] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
				else
				begin
					map[55:52] <= map[63:60];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
			end
			else if (map[63:60] > 0 && map[59:56] == 0 && map[55:52] > 0 && map[51:48] == 0)
			begin
				if (map[55:52] == map[63:60])
				begin
					map[51:48] <= (map[63:60] + 1);
					map[63:60] <= 0;
					map[55:52] <= 1;
				end
				else
				begin
					map[51:48] <= map[55:52];
					map[55:52] <= map[63:60];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
			end
			else if (map[63:60] > 0 && map[59:56] > 0 && map[55:52] == 0 && map[51:48] == 0)
			begin
				if (map[59:56] == map[63:60])
				begin
					map[51:48] <= (map[63:60] + 1);
					map[63:60] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
					   	map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
				else
				begin
					map[51:48] <= map[59:56];
					map[55:52] <= map[63:60];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
					map[63:60] <= 0;
				end
			end
			else if (map[63:60] > 0 && map[59:56] > 0 && map[55:52] > 0 && map[51:48] == 0)
			begin
				if (map[55:52] == map[59:56])
				begin
					map[51:48] <= (map[55:52] + 1);
					map[55:52] <= map[63:60];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
					map[59:56] <= 0;
				end
				else
				if (map[63:60] == map[59:56])
				begin
					map[51:48] <= map[55:52];
					map[55:52] <= (map[59:56] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
					map[59:56] <= 0;
				end
				else
				begin
					map[51:48] <= map[55:52];
					map[55:52] <= map[59:56];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
					map[59:56] <= map[63:60];
				end
			end
			else if (map[63:60] > 0 && map[59:56] == 0 && map[55:52] > 0 && map[51:48] > 0)
			begin
				if (map[55:52] == map[51:48])
				begin
					map[51:48] <= (map[51:48] + 1);
					map[55:52] <= map[63:60];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
					    map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
					map[63:60] <= 0;
				end
				else
				if (map[63:60] == map[55:52])
				begin
					map[55:52] <= (map[55:52] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
				else
				begin
					map[59:56] <= map[63:60];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
			end
			else if (map[63:60] > 0 && map[59:56] > 0 && map[55:52] == 0 && map[51:48] > 0)
			begin
				if (map[59:56] == map[51:48])
				begin
					map[51:48] <= (map[51:48] + 1);
					map[55:52] <= map[63:60];
					map[59:56] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
				else
				if (map[63:60] == map[59:56])
				begin
					map[55:52] <= (map[59:56] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
					map[59:56] <= 0;
				end
				else
				begin
					map[55:52] <= map[59:56];
					map[59:56] <= map[63:60];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
			end
			else if (map[63:60] > 0 && map[59:56] > 0 && map[55:52] > 0 && map[51:48] > 0)
			begin
				if (map[55:52] == map[51:48])
				begin
					map[51:48] <= (map[51:48] + 1);
					if (map[63:60] == map[59:56])
					begin
						map[55:52] <= (map[59:56] + 1);
						if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
						begin
							map[63:60] <= 1;
						end
						else
						begin
							map[63:60] <= 0;
						end
						map[59:56] <= 0;
					end
					else
					begin
						map[55:52] <= map[59:56];
						if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
						begin
							map[63:60] <= 1;
						end
						else
						begin
							map[63:60] <= 0;
						end
						map[59:56] <= map[63:60];
					end
				end
				else
				if (map[59:56] == map[55:52])
				begin
					map[55:52] <= (map[55:52] + 1);
					map[59:56] <= map[63:60];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
				else
				if (map[63:60] == map[59:56])
				begin
					map[59:56] <= (map[59:56] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[63:60] <= 1;
					end
					else
					begin
						map[63:60] <= 0;
					end
				end
			end
			else if (map[63:60] == 0 && map[59:56] > 0 && map[55:52] == 0 && map[51:48] == 0)
			begin
				map[51:48] <= map[59:56];
				if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
				begin
					map[59:56] <= 1;
				end
				else
				begin
					map[59:56] <= 0;
				end
			end
			else if (map[63:60] == 0 && map[59:56] == 0 && map[55:52] > 0 && map[51:48] == 0)
			begin
				map[51:48] <= map[55:52];
				map[55:52] <= 1;
			end
			else if (map[63:60] == 0 && map[59:56] == 0 && map[55:52] == 0 && map[51:48] > 0)
			begin
			end
			else if (map[63:60] == 0 && map[59:56] > 0 && map[55:52] == 0 && map[51:48] > 0)
			begin
				if (map[51:48] == map[59:56])
				begin
					map[51:48] <= (map[51:48] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
				else
				begin
					map[55:52] <= map[59:56];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
			end
			else if (map[63:60] == 0 && map[59:56] == 0 && map[55:52] > 0 && map[51:48] > 0)
			begin
				if (map[55:52] == map[51:48])
				begin
					map[51:48] <= (map[51:48] + 1);
					map[55:52] <= 1;
				end
			end
			else if (map[63:60] == 0 && map[59:56] > 0 && map[55:52] > 0 && map[51:48] == 0)
			begin
				if (map[59:56] == map[55:52])
				begin
					map[51:48] <= (map[55:52] + 1);
					map[55:52] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
				else
				begin
					map[51:48] <= map[55:52];
					map[55:52] <= map[59:56];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
			end
			else if (map[63:60] == 0 && map[59:56] > 0 && map[55:52] > 0 && map[51:48] > 0)
			begin
				if (map[51:48] == map[55:52])
				begin
					map[51:48] <= (map[55:52] + 1);
					map[55:52] <= map[59:56];
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
				else
				if (map[55:52] == map[59:56])
				begin
					map[55:52] <= (map[55:52] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[15:12] != map[11:8] && map[11:8] != map[7:4] && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] == 0) || 
						(map[15:12] == 0 && map[11:8] > 0 && map[7:4] > 0 && map[3:0] > 0 && map[11:8] != map[7:4] && map[7:4] != map[3:0]) ||
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] > 0 && map[3:0] > 0 && map[7:4] != map[3:0]) || 
						(map[15:12] == 0 && map[11:8] == 0 && map[7:4] == 0 && map[3:0] > 0)
					)
					&& 
					(
						(map[31:28] > 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[31:28] != map[27:24] && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] == 0) || 
						(map[31:28] == 0 && map[27:24] > 0 && map[23:20] > 0 && map[19:16] > 0 && map[27:24] != map[23:20] && map[23:20] != map[19:16]) ||
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] > 0 && map[19:16] > 0 && map[23:20] != map[19:16]) || 
						(map[31:28] == 0 && map[27:24] == 0 && map[23:20] == 0 && map[19:16] > 0)
					)
					&& 
					(	
						(map[47:44] > 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[47:44] != map[43:40] && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] == 0) || 
						(map[47:44] == 0 && map[43:40] > 0 && map[39:36] > 0 && map[35:32] > 0 && map[43:40] != map[39:36] && map[39:36] != map[35:32]) ||
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] > 0 && map[35:32] > 0 && map[39:36] != map[35:32]) || 
						(map[47:44] == 0 && map[43:40] == 0 && map[39:36] == 0 && map[35:32] > 0)
					)
				)
					begin
						map[59:56] <= 1;
					end
					else
					begin
						map[59:56] <= 0;
					end
				end
			end
			else if (map[63:60] == 0 && map[59:56] == 0 && map[55:52] == 0 && map[51:48] == 0)
			begin
			end
		end
		else
		if (down == 1)
		begin
			/*Down*/
			/*First line*/
			if (map[15:12] > 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0)
			begin
				map[63:60] <= map[15:12];
				map[15:12] <= 1;
			end
			else if (map[15:12] > 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
			begin
				if (map[63:60] == map[15:12])
				begin
					map[63:60] <= (map[15:12] + 1);
					map[15:12] <= 1;
				end
				else
				begin
					map[47:44] <= map[15:12];
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] > 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] == 0)
			begin
				if (map[47:44] == map[15:12])
				begin
					map[63:60] <= (map[15:12] + 1);
					map[15:12] <= 0;
					map[47:44] <= 1;
				end
				else
				begin
					map[63:60] <= map[47:44];
					map[47:44] <= map[15:12];
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] > 0 && map[31:28] > 0 && map[47:44] == 0 && map[63:60] == 0)
			begin
				if (map[31:28] == map[15:12])
				begin
					map[63:60] <= (map[15:12] + 1);
					map[15:12] <= 0;
					map[31:28] <= 1;
				end
				else
				begin
					map[63:60] <= map[31:28];
					map[47:44] <= map[15:12];
					map[31:28] <= 1;
					map[15:12] <= 0;
				end
			end
			else if (map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] == 0)
			begin
				if (map[47:44] == map[31:28])
				begin
					map[63:60] <= (map[47:44] + 1);
					map[47:44] <= map[15:12];
					map[15:12] <= 1;
					map[31:28] <= 0;
				end
				else
				if (map[15:12] == map[31:28])
				begin
					map[63:60] <= map[47:44];
					map[47:44] <= (map[31:28] + 1);
					map[15:12] <= 1;
					map[31:28] <= 0;
				end
				else
				begin
					map[63:60] <= map[47:44];
					map[47:44] <= map[31:28];
					map[15:12] <= 1;
					map[31:28] <= map[15:12];
				end
			end
			else if (map[15:12] > 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0)
			begin
				if (map[47:44] == map[63:60])
				begin
					map[63:60] <= (map[63:60] + 1);
					map[47:44] <= map[15:12];
					map[31:28] <= 1;
					map[15:12] <= 0;
				end
				else
				if (map[15:12] == map[47:44])
				begin
					map[47:44] <= (map[47:44] + 1);
					map[15:12] <= 1;
				end
				else
				begin
					map[31:28] <= map[15:12];
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] > 0 && map[31:28] > 0 && map[47:44] == 0 && map[63:60] > 0)
			begin
				if (map[31:28] == map[63:60])
				begin
					map[63:60] <= (map[63:60] + 1);
					map[47:44] <= map[15:12];
					map[31:28] <= 0;
					map[15:12] <= 1;
				end
				else
				if (map[15:12] == map[31:28])
				begin
					map[47:44] <= (map[31:28] + 1);
					map[15:12] <= 1;
					map[31:28] <= 0;
				end
				else
				begin
					map[47:44] <= map[31:28];
					map[31:28] <= map[15:12];
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0)
			begin
				if (map[47:44] == map[63:60])
				begin
					map[63:60] <= (map[63:60] + 1);
					if (map[15:12] == map[31:28])
					begin
						map[47:44] <= (map[31:28] + 1);
						map[15:12] <= 1;
						map[31:28] <= 0;
					end
					else
					begin
						map[47:44] <= map[31:28];
						map[15:12] <= 1;
						map[31:28] <= map[15:12];
					end
				end
				else
				if (map[31:28] == map[47:44])
				begin
					map[47:44] <= (map[47:44] + 1);
					map[31:28] <= map[15:12];
					map[15:12] <= 1;
				end
				else
				if (map[15:12] == map[31:28])
				begin
					map[31:28] <= (map[31:28] + 1);
					map[15:12] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[31:28] > 0 && map[47:44] == 0 && map[63:60] == 0)
			begin
				map[63:60] <= map[31:28];
				map[31:28] <= 1;
			end
			else if (map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] == 0)
			begin
				map[63:60] <= map[47:44];
				map[47:44] <= 1;
			end
			else if (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
			begin
			end
			else if (map[15:12] == 0 && map[31:28] > 0 && map[47:44] == 0 && map[63:60] > 0)
			begin
				if (map[63:60] == map[31:28])
				begin
					map[63:60] <= (map[63:60] + 1);
					map[31:28] <= 1;
				end
				else
				begin
					map[47:44] <= map[31:28];
					map[31:28] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0)
			begin
				if (map[47:44] == map[63:60])
				begin
					map[63:60] <= (map[63:60] + 1);
					map[47:44] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] == 0)
			begin
				if (map[31:28] == map[47:44])
				begin
					map[63:60] <= (map[47:44] + 1);
					map[47:44] <= 0;
					map[31:28] <= 1;
				end
				else
				begin
					map[63:60] <= map[47:44];
					map[47:44] <= map[31:28];
					map[31:28] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0)
			begin
				if (map[63:60] == map[47:44])
				begin
					map[63:60] <= (map[47:44] + 1);
					map[47:44] <= map[31:28];
					map[31:28] <= 1;
				end
				else
				if (map[47:44] == map[31:28])
				begin
					map[47:44] <= (map[47:44] + 1);
					map[31:28] <= 1;
				end
			end
			else if (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0)
			begin
			end
			
			/*Second line*/			
			
			if (map[11:8] > 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0)
			begin
				map[59:56] <= map[11:8];
				if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
				begin
					map[11:8] <= 1;
				end
				else
				begin
					map[11:8] <= 0;
				end
			end
			else if (map[11:8] > 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
			begin
				if (map[59:56] == map[11:8])
				begin
					map[59:56] <= (map[11:8] + 1);
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
				else
				begin
					map[43:40] <= map[11:8];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
			end
			else if (map[11:8] > 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] == 0)
			begin
				if (map[43:40] == map[11:8])
				begin
					map[59:56] <= (map[11:8] + 1);
					map[11:8] <= 0;
					map[43:40] <= 1;
				end
				else
				begin
					map[59:56] <= map[43:40];
					map[43:40] <= map[11:8];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
			end
			else if (map[11:8] > 0 && map[27:24] > 0 && map[43:40] == 0 && map[59:56] == 0)
			begin
				if (map[27:24] == map[11:8])
				begin
					map[59:56] <= (map[11:8] + 1);
					map[11:8] <= 0;
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
					   	map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
				else
				begin
					map[59:56] <= map[27:24];
					map[43:40] <= map[11:8];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
					map[11:8] <= 0;
				end
			end
			else if (map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] == 0)
			begin
				if (map[43:40] == map[27:24])
				begin
					map[59:56] <= (map[43:40] + 1);
					map[43:40] <= map[11:8];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
					map[27:24] <= 0;
				end
				else
				if (map[11:8] == map[27:24])
				begin
					map[59:56] <= map[43:40];
					map[43:40] <= (map[27:24] + 1);
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
					map[27:24] <= 0;
				end
				else
				begin
					map[59:56] <= map[43:40];
					map[43:40] <= map[27:24];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
					map[27:24] <= map[11:8];
				end
			end
			else if (map[11:8] > 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0)
			begin
				if (map[43:40] == map[59:56])
				begin
					map[59:56] <= (map[59:56] + 1);
					map[43:40] <= map[11:8];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
					    map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
					map[11:8] <= 0;
				end
				else
				if (map[11:8] == map[43:40])
				begin
					map[43:40] <= (map[43:40] + 1);
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
				else
				begin
					map[27:24] <= map[11:8];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
			end
			else if (map[11:8] > 0 && map[27:24] > 0 && map[43:40] == 0 && map[59:56] > 0)
			begin
				if (map[27:24] == map[59:56])
				begin
					map[59:56] <= (map[59:56] + 1);
					map[43:40] <= map[11:8];
					map[27:24] <= 0;
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
				else
				if (map[11:8] == map[27:24])
				begin
					map[43:40] <= (map[27:24] + 1);
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
					map[27:24] <= 0;
				end
				else
				begin
					map[43:40] <= map[27:24];
					map[27:24] <= map[11:8];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
			end
			else if (map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0)
			begin
				if (map[43:40] == map[59:56])
				begin
					map[59:56] <= (map[59:56] + 1);
					if (map[11:8] == map[27:24])
					begin
						map[43:40] <= (map[27:24] + 1);
						if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
						begin
							map[11:8] <= 1;
						end
						else
						begin
							map[11:8] <= 0;
						end
						map[27:24] <= 0;
					end
					else
					begin
						map[43:40] <= map[27:24];
						if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
						begin
							map[11:8] <= 1;
						end
						else
						begin
							map[11:8] <= 0;
						end
						map[27:24] <= map[11:8];
					end
				end
				else
				if (map[27:24] == map[43:40])
				begin
					map[43:40] <= (map[43:40] + 1);
					map[27:24] <= map[11:8];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
				else
				if (map[11:8] == map[27:24])
				begin
					map[27:24] <= (map[27:24] + 1);
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[11:8] <= 1;
					end
					else
					begin
						map[11:8] <= 0;
					end
				end
			end
			else if (map[11:8] == 0 && map[27:24] > 0 && map[43:40] == 0 && map[59:56] == 0)
			begin
				map[59:56] <= map[27:24];
				if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
				begin
					map[27:24] <= 1;
				end
				else
				begin
					map[27:24] <= 0;
				end
			end
			else if (map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] == 0)
			begin
				map[59:56] <= map[43:40];
				map[43:40] <= 1;
			end
			else if (map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
			begin
			end
			else if (map[11:8] == 0 && map[27:24] > 0 && map[43:40] == 0 && map[59:56] > 0)
			begin
				if (map[59:56] == map[27:24])
				begin
					map[59:56] <= (map[59:56] + 1);
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
				else
				begin
					map[43:40] <= map[27:24];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
			end
			else if (map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0)
			begin
				if (map[43:40] == map[59:56])
				begin
					map[59:56] <= (map[59:56] + 1);
					map[43:40] <= 1;
				end
			end
			else if (map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] == 0)
			begin
				if (map[27:24] == map[43:40])
				begin
					map[59:56] <= (map[43:40] + 1);
					map[43:40] <= 0;
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
				else
				begin
					map[59:56] <= map[43:40];
					map[43:40] <= map[27:24];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
			end
			else if (map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0)
			begin
				if (map[59:56] == map[43:40])
				begin
					map[59:56] <= (map[43:40] + 1);
					map[43:40] <= map[27:24];
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
				else
				if (map[43:40] == map[27:24])
				begin
					map[43:40] <= (map[43:40] + 1);
					if ((map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0
				&& map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || (map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
				(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || (map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0))
					begin
						map[27:24] <= 1;
					end
					else
					begin
						map[27:24] <= 0;
					end
				end
			end
			else if (map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0)
			begin
			end

			/*Third line*/			
			
			if (map[7:4] > 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0)
			begin
				map[55:52] <= map[7:4];
				if 
				( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
				begin
					map[7:4] <= 1;
				end
				else
				begin
					map[7:4] <= 0;
				end
			end
			else if (map[7:4] > 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
			begin
				if (map[55:52] == map[7:4])
				begin
					map[55:52] <= (map[7:4] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
				else
				begin
					map[39:36] <= map[7:4];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
			end
			else if (map[7:4] > 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] == 0)
			begin
				if (map[39:36] == map[7:4])
				begin
					map[55:52] <= (map[7:4] + 1);
					map[7:4] <= 0;
					map[39:36] <= 1;
				end
				else
				begin
					map[55:52] <= map[39:36];
					map[39:36] <= map[7:4];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
			end
			else if (map[7:4] > 0 && map[23:20] > 0 && map[39:36] == 0 && map[55:52] == 0)
			begin
				if (map[23:20] == map[7:4])
				begin
					map[55:52] <= (map[7:4] + 1);
					map[7:4] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
					   	map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
				else
				begin
					map[55:52] <= map[23:20];
					map[39:36] <= map[7:4];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
					map[7:4] <= 0;
				end
			end
			else if (map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] == 0)
			begin
				if (map[39:36] == map[23:20])
				begin
					map[55:52] <= (map[39:36] + 1);
					map[39:36] <= map[7:4];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
					map[23:20] <= 0;
				end
				else
				if (map[7:4] == map[23:20])
				begin
					map[55:52] <= map[39:36];
					map[39:36] <= (map[23:20] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
					map[23:20] <= 0;
				end
				else
				begin
					map[55:52] <= map[39:36];
					map[39:36] <= map[23:20];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
					map[23:20] <= map[7:4];
				end
			end
			else if (map[7:4] > 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0)
			begin
				if (map[39:36] == map[55:52])
				begin
					map[55:52] <= (map[55:52] + 1);
					map[39:36] <= map[7:4];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
					    map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
					map[7:4] <= 0;
				end
				else
				if (map[7:4] == map[39:36])
				begin
					map[39:36] <= (map[39:36] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
				else
				begin
					map[23:20] <= map[7:4];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
			end
			else if (map[7:4] > 0 && map[23:20] > 0 && map[39:36] == 0 && map[55:52] > 0)
			begin
				if (map[23:20] == map[55:52])
				begin
					map[55:52] <= (map[55:52] + 1);
					map[39:36] <= map[7:4];
					map[23:20] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
				else
				if (map[7:4] == map[23:20])
				begin
					map[39:36] <= (map[23:20] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
					map[23:20] <= 0;
				end
				else
				begin
					map[39:36] <= map[23:20];
					map[23:20] <= map[7:4];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
			end
			else if (map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0)
			begin
				if (map[39:36] == map[55:52])
				begin
					map[55:52] <= (map[55:52] + 1);
					if (map[7:4] == map[23:20])
					begin
						map[39:36] <= (map[23:20] + 1);
						if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
						begin
							map[7:4] <= 1;
						end
						else
						begin
							map[7:4] <= 0;
						end
						map[23:20] <= 0;
					end
					else
					begin
						map[39:36] <= map[23:20];
						if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
						begin
							map[7:4] <= 1;
						end
						else
						begin
							map[7:4] <= 0;
						end
						map[23:20] <= map[7:4];
					end
				end
				else
				if (map[23:20] == map[39:36])
				begin
					map[39:36] <= (map[39:36] + 1);
					map[23:20] <= map[7:4];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
				else
				if (map[7:4] == map[23:20])
				begin
					map[23:20] <= (map[23:20] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[7:4] <= 1;
					end
					else
					begin
						map[7:4] <= 0;
					end
				end
			end
			else if (map[7:4] == 0 && map[23:20] > 0 && map[39:36] == 0 && map[55:52] == 0)
			begin
				map[55:52] <= map[23:20];
				if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
				begin
					map[23:20] <= 1;
				end
				else
				begin
					map[23:20] <= 0;
				end
			end
			else if (map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] == 0)
			begin
				map[55:52] <= map[39:36];
				map[39:36] <= 1;
			end
			else if (map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
			begin
			end
			else if (map[7:4] == 0 && map[23:20] > 0 && map[39:36] == 0 && map[55:52] > 0)
			begin
				if (map[55:52] == map[23:20])
				begin
					map[55:52] <= (map[55:52] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
				else
				begin
					map[39:36] <= map[23:20];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
			end
			else if (map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0)
			begin
				if (map[39:36] == map[55:52])
				begin
					map[55:52] <= (map[55:52] + 1);
					map[39:36] <= 1;
				end
			end
			else if (map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] == 0)
			begin
				if (map[23:20] == map[39:36])
				begin
					map[55:52] <= (map[39:36] + 1);
					map[39:36] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
				else
				begin
					map[55:52] <= map[39:36];
					map[39:36] <= map[23:20];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
			end
			else if (map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0)
			begin
				if (map[55:52] == map[39:36])
				begin
					map[55:52] <= (map[39:36] + 1);
					map[39:36] <= map[23:20];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
				else
				if (map[39:36] == map[23:20])
				begin
					map[39:36] <= (map[39:36] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
				)	
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
			end
			else if (map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0)
			begin
			end

			/*Forth line*/			
			
			if (map[3:0] > 0 && map[19:16] == 0 && map[35:32] == 0 && map[51:48] == 0)
			begin
				map[51:48] <= map[3:0];
				if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
				begin
					map[3:0] <= 1;
				end
				else
				begin
					map[3:0] <= 0;
				end
			end
			else if (map[3:0] > 0 && map[19:16] == 0 && map[35:32] == 0 && map[51:48] > 0)
			begin
				if (map[51:48] == map[3:0])
				begin
					map[51:48] <= (map[3:0] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
				else
				begin
					map[35:32] <= map[3:0];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
			end
			else if (map[3:0] > 0 && map[19:16] == 0 && map[35:32] > 0 && map[51:48] == 0)
			begin
				if (map[35:32] == map[3:0])
				begin
					map[51:48] <= (map[3:0] + 1);
					map[3:0] <= 0;
					map[35:32] <= 1;
				end
				else
				begin
					map[51:48] <= map[35:32];
					map[35:32] <= map[3:0];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
			end
			else if (map[3:0] > 0 && map[19:16] > 0 && map[35:32] == 0 && map[51:48] == 0)
			begin
				if (map[19:16] == map[3:0])
				begin
					map[51:48] <= (map[3:0] + 1);
					map[3:0] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
					   	map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
				else
				begin
					map[51:48] <= map[19:16];
					map[35:32] <= map[3:0];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
					map[3:0] <= 0;
				end
			end
			else if (map[3:0] > 0 && map[19:16] > 0 && map[35:32] > 0 && map[51:48] == 0)
			begin
				if (map[35:32] == map[19:16])
				begin
					map[51:48] <= (map[35:32] + 1);
					map[35:32] <= map[3:0];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
					map[19:16] <= 0;
				end
				else
				if (map[3:0] == map[19:16])
				begin
					map[51:48] <= map[35:32];
					map[35:32] <= (map[19:16] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
					map[19:16] <= 0;
				end
				else
				begin
					map[51:48] <= map[35:32];
					map[35:32] <= map[19:16];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
					map[19:16] <= map[3:0];
				end
			end
			else if (map[3:0] > 0 && map[19:16] == 0 && map[35:32] > 0 && map[51:48] > 0)
			begin
				if (map[35:32] == map[51:48])
				begin
					map[51:48] <= (map[51:48] + 1);
					map[35:32] <= map[3:0];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
					    map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
					map[3:0] <= 0;
				end
				else
				if (map[3:0] == map[35:32])
				begin
					map[35:32] <= (map[35:32] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
				else
				begin
					map[19:16] <= map[3:0];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
			end
			else if (map[3:0] > 0 && map[19:16] > 0 && map[35:32] == 0 && map[51:48] > 0)
			begin
				if (map[19:16] == map[51:48])
				begin
					map[51:48] <= (map[51:48] + 1);
					map[35:32] <= map[3:0];
					map[19:16] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
				else
				if (map[3:0] == map[19:16])
				begin
					map[35:32] <= (map[19:16] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
					map[19:16] <= 0;
				end
				else
				begin
					map[35:32] <= map[19:16];
					map[19:16] <= map[3:0];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
			end
			else if (map[3:0] > 0 && map[19:16] > 0 && map[35:32] > 0 && map[51:48] > 0)
			begin
				if (map[35:32] == map[51:48])
				begin
					map[51:48] <= (map[51:48] + 1);
					if (map[3:0] == map[19:16])
					begin
						map[35:32] <= (map[19:16] + 1);
						if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
						begin
							map[3:0] <= 1;
						end
						else
						begin
							map[3:0] <= 0;
						end
						map[19:16] <= 0;
					end
					else
					begin
						map[35:32] <= map[19:16];
						if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
						begin
							map[3:0] <= 1;
						end
						else
						begin
							map[3:0] <= 0;
						end
						map[19:16] <= map[3:0];
					end
				end
				else
				if (map[19:16] == map[35:32])
				begin
					map[35:32] <= (map[35:32] + 1);
					map[19:16] <= map[3:0];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
				else
				if (map[3:0] == map[19:16])
				begin
					map[19:16] <= (map[19:16] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[3:0] <= 1;
					end
					else
					begin
						map[3:0] <= 0;
					end
				end
			end
			else if (map[3:0] == 0 && map[19:16] > 0 && map[35:32] == 0 && map[51:48] == 0)
			begin
				map[51:48] <= map[19:16];
				if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
				begin
					map[19:16] <= 1;
				end
				else
				begin
					map[19:16] <= 0;
				end
			end
			else if (map[3:0] == 0 && map[19:16] == 0 && map[35:32] > 0 && map[51:48] == 0)
			begin
				map[51:48] <= map[35:32];
				map[35:32] <= 1;
			end
			else if (map[3:0] == 0 && map[19:16] == 0 && map[35:32] == 0 && map[51:48] > 0)
			begin
			end
			else if (map[3:0] == 0 && map[19:16] > 0 && map[35:32] == 0 && map[51:48] > 0)
			begin
				if (map[51:48] == map[19:16])
				begin
					map[51:48] <= (map[51:48] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
				else
				begin
					map[35:32] <= map[19:16];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
			end
			else if (map[3:0] == 0 && map[19:16] == 0 && map[35:32] > 0 && map[51:48] > 0)
			begin
				if (map[35:32] == map[51:48])
				begin
					map[51:48] <= (map[51:48] + 1);
					map[35:32] <= 1;
				end
			end
			else if (map[3:0] == 0 && map[19:16] > 0 && map[35:32] > 0 && map[51:48] == 0)
			begin
				if (map[19:16] == map[35:32])
				begin
					map[51:48] <= (map[35:32] + 1);
					map[35:32] <= 0;
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
				else
				begin
					map[51:48] <= map[35:32];
					map[35:32] <= map[19:16];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
			end
			else if (map[3:0] == 0 && map[19:16] > 0 && map[35:32] > 0 && map[51:48] > 0)
			begin
				if (map[51:48] == map[35:32])
				begin
					map[51:48] <= (map[35:32] + 1);
					map[35:32] <= map[19:16];
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
				else
				if (map[35:32] == map[19:16])
				begin
					map[35:32] <= (map[35:32] + 1);
					if ( 
					( 
						(map[15:12] > 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[15:12] != map[31:28] && map[31:28] != map[47:44] && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] == 0) || 
						(map[15:12] == 0 && map[31:28] > 0 && map[47:44] > 0 && map[63:60] > 0 && map[31:28] != map[47:44] && map[47:44] != map[63:60]) ||
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] > 0 && map[63:60] > 0 && map[47:44] != map[63:60]) || 
						(map[15:12] == 0 && map[31:28] == 0 && map[47:44] == 0 && map[63:60] > 0)
					)
					&& 
					(
						(map[11:8] > 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[11:8] != map[27:24] && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] == 0) || 
						(map[11:8] == 0 && map[27:24] > 0 && map[43:40] > 0 && map[59:56] > 0 && map[27:24] != map[43:40] && map[43:40] != map[59:56]) ||
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] > 0 && map[59:56] > 0 && map[43:40] != map[59:56]) || 
						(map[11:8] == 0 && map[27:24] == 0 && map[43:40] == 0 && map[59:56] > 0)
					)
					&& 
					(	
						(map[7:4] > 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[7:4] != map[23:20] && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] == 0) || 
						(map[7:4] == 0 && map[23:20] > 0 && map[39:36] > 0 && map[55:52] > 0 && map[23:20] != map[39:36] && map[39:36] != map[55:52]) ||
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] > 0 && map[55:52] > 0 && map[39:36] != map[55:52]) || 
						(map[7:4] == 0 && map[23:20] == 0 && map[39:36] == 0 && map[55:52] > 0)
					)
				)
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
			end
			else if (map[3:0] == 0 && map[19:16] == 0 && map[35:32] == 0 && map[51:48] == 0)
			begin
			end
		end
		else
		if (right == 1)
		begin
			/*Right*/
			/*First line*/
			if (map[3:0] > 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0)
			begin
				map[15:12] <= map[3:0];
				map[3:0] <= 1;
			end
			else if (map[3:0] > 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
			begin
				if (map[15:12] == map[3:0])
				begin
					map[15:12] <= (map[3:0] + 1);
					map[3:0] <= 1;
				end
				else
				begin
					map[11:8] <= map[3:0];
					map[3:0] <= 1;
				end
			end
			else if (map[3:0] > 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] == 0)
			begin
				if (map[11:8] == map[3:0])
				begin
					map[15:12] <= (map[3:0] + 1);
					map[3:0] <= 0;
					map[11:8] <= 1;
				end
				else
				begin
					map[15:12] <= map[11:8];
					map[11:8] <= map[3:0];
					map[3:0] <= 1;
				end
			end
			else if (map[3:0] > 0 && map[7:4] > 0 && map[11:8] == 0 && map[15:12] == 0)
			begin
				if (map[7:4] == map[3:0])
				begin
					map[15:12] <= (map[3:0] + 1);
					map[3:0] <= 0;
					map[7:4] <= 1;
				end
				else
				begin
					map[15:12] <= map[7:4];
					map[11:8] <= map[3:0];
					map[7:4] <= 1;
					map[3:0] <= 0;
				end
			end
			else if (map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] == 0)
			begin
				if (map[11:8] == map[7:4])
				begin
					map[15:12] <= (map[11:8] + 1);
					map[11:8] <= map[3:0];
					map[3:0] <= 1;
					map[7:4] <= 0;
				end
				else
				if (map[3:0] == map[7:4])
				begin
					map[15:12] <= map[11:8];
					map[11:8] <= (map[7:4] + 1);
					map[3:0] <= 1;
					map[7:4] <= 0;
				end
				else
				begin
					map[15:12] <= map[11:8];
					map[11:8] <= map[7:4];
					map[3:0] <= 1;
					map[7:4] <= map[3:0];
				end
			end
			else if (map[3:0] > 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0)
			begin
				if (map[11:8] == map[15:12])
				begin
					map[15:12] <= (map[15:12] + 1);
					map[11:8] <= map[3:0];
					map[7:4] <= 1;
					map[3:0] <= 0;
				end
				else
				if (map[3:0] == map[11:8])
				begin
					map[11:8] <= (map[11:8] + 1);
					map[3:0] <= 1;
				end
				else
				begin
					map[7:4] <= map[3:0];
					map[3:0] <= 1;
				end
			end
			else if (map[3:0] > 0 && map[7:4] > 0 && map[11:8] == 0 && map[15:12] > 0)
			begin
				if (map[7:4] == map[15:12])
				begin
					map[15:12] <= (map[15:12] + 1);
					map[11:8] <= map[3:0];
					map[7:4] <= 0;
					map[3:0] <= 1;
				end
				else
				if (map[3:0] == map[7:4])
				begin
					map[11:8] <= (map[7:4] + 1);
					map[3:0] <= 1;
					map[7:4] <= 0;
				end
				else
				begin
					map[11:8] <= map[7:4];
					map[7:4] <= map[3:0];
					map[3:0] <= 1;
				end
			end
			else if (map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0)
			begin
				if (map[11:8] == map[15:12])
				begin
					map[15:12] <= (map[15:12] + 1);
					if (map[3:0] == map[7:4])
					begin
						map[11:8] <= (map[7:4] + 1);
						map[3:0] <= 1;
						map[7:4] <= 0;
					end
					else
					begin
						map[11:8] <= map[7:4];
						map[3:0] <= 1;
						map[7:4] <= map[3:0];
					end
				end
				else
				if (map[7:4] == map[11:8])
				begin
					map[11:8] <= (map[11:8] + 1);
					map[7:4] <= map[3:0];
					map[3:0] <= 1;
				end
				else
				if (map[3:0] == map[7:4])
				begin
					map[7:4] <= (map[7:4] + 1);
					map[3:0] <= 1;
				end
			end
			else if (map[3:0] == 0 && map[7:4] > 0 && map[11:8] == 0 && map[15:12] == 0)
			begin
				map[15:12] <= map[7:4];
				map[7:4] <= 1;
			end
			else if (map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] == 0)
			begin
				map[15:12] <= map[11:8];
				map[11:8] <= 1;
			end
			else if (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
			begin
			end
			else if (map[3:0] == 0 && map[7:4] > 0 && map[11:8] == 0 && map[15:12] > 0)
			begin
				if (map[15:12] == map[7:4])
				begin
					map[15:12] <= (map[15:12] + 1);
					map[7:4] <= 1;
				end
				else
				begin
					map[11:8] <= map[7:4];
					map[7:4] <= 1;
				end
			end
			else if (map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0)
			begin
				if (map[11:8] == map[15:12])
				begin
					map[15:12] <= (map[15:12] + 1);
					map[11:8] <= 1;
				end
			end
			else if (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] == 0)
			begin
				if (map[7:4] == map[11:8])
				begin
					map[15:12] <= (map[11:8] + 1);
					map[11:8] <= 0;
					map[7:4] <= 1;
				end
				else
				begin
					map[15:12] <= map[11:8];
					map[11:8] <= map[7:4];
					map[7:4] <= 1;
				end
			end
			else if (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0)
			begin
				if (map[15:12] == map[11:8])
				begin
					map[15:12] <= (map[11:8] + 1);
					map[11:8] <= map[7:4];
					map[7:4] <= 1;
				end
				else
				if (map[11:8] == map[7:4])
				begin
					map[11:8] <= (map[11:8] + 1);
					map[7:4] <= 1;
				end
			end
			else if (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0)
			begin
			end
			
			/*Second line*/			
			
			if (map[19:16] > 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0)
			begin
				map[31:28] <= map[19:16];
				if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
				begin
					map[19:16] <= 1;
				end
				else
				begin
					map[19:16] <= 0;
				end
			end
			else if (map[19:16] > 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
			begin
				if (map[31:28] == map[19:16])
				begin
					map[31:28] <= (map[19:16] + 1);
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
				else
				begin
					map[27:24] <= map[19:16];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
			end
			else if (map[19:16] > 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] == 0)
			begin
				if (map[27:24] == map[19:16])
				begin
					map[31:28] <= (map[19:16] + 1);
					map[19:16] <= 0;
					map[27:24] <= 1;
				end
				else
				begin
					map[31:28] <= map[27:24];
					map[27:24] <= map[19:16];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
			end
			else if (map[19:16] > 0 && map[23:20] > 0 && map[27:24] == 0 && map[31:28] == 0)
			begin
				if (map[23:20] == map[19:16])
				begin
					map[31:28] <= (map[19:16] + 1);
					map[19:16] <= 0;
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
					   	map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
				else
				begin
					map[31:28] <= map[23:20];
					map[27:24] <= map[19:16];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
					map[19:16] <= 0;
				end
			end
			else if (map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] == 0)
			begin
				if (map[27:24] == map[23:20])
				begin
					map[31:28] <= (map[27:24] + 1);
					map[27:24] <= map[19:16];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
					map[23:20] <= 0;
				end
				else
				if (map[19:16] == map[23:20])
				begin
					map[31:28] <= map[27:24];
					map[27:24] <= (map[23:20] + 1);
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
					map[23:20] <= 0;
				end
				else
				begin
					map[31:28] <= map[27:24];
					map[27:24] <= map[23:20];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
					map[23:20] <= map[19:16];
				end
			end
			else if (map[19:16] > 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0)
			begin
				if (map[27:24] == map[31:28])
				begin
					map[31:28] <= (map[31:28] + 1);
					map[27:24] <= map[19:16];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
					    map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
					map[19:16] <= 0;
				end
				else
				if (map[19:16] == map[27:24])
				begin
					map[27:24] <= (map[27:24] + 1);
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
				else
				begin
					map[23:20] <= map[19:16];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
			end
			else if (map[19:16] > 0 && map[23:20] > 0 && map[27:24] == 0 && map[31:28] > 0)
			begin
				if (map[23:20] == map[31:28])
				begin
					map[31:28] <= (map[31:28] + 1);
					map[27:24] <= map[19:16];
					map[23:20] <= 0;
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
				else
				if (map[19:16] == map[23:20])
				begin
					map[27:24] <= (map[23:20] + 1);
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
					map[23:20] <= 0;
				end
				else
				begin
					map[27:24] <= map[23:20];
					map[23:20] <= map[19:16];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
			end
			else if (map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0)
			begin
				if (map[27:24] == map[31:28])
				begin
					map[31:28] <= (map[31:28] + 1);
					if (map[19:16] == map[23:20])
					begin
						map[27:24] <= (map[23:20] + 1);
						if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
						begin
							map[19:16] <= 1;
						end
						else
						begin
							map[19:16] <= 0;
						end
						map[23:20] <= 0;
					end
					else
					begin
						map[27:24] <= map[23:20];
						if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
						begin
							map[19:16] <= 1;
						end
						else
						begin
							map[19:16] <= 0;
						end
						map[23:20] <= map[19:16];
					end
				end
				else
				if (map[23:20] == map[27:24])
				begin
					map[27:24] <= (map[27:24] + 1);
					map[23:20] <= map[19:16];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
				else
				if (map[19:16] == map[23:20])
				begin
					map[23:20] <= (map[23:20] + 1);
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[19:16] <= 1;
					end
					else
					begin
						map[19:16] <= 0;
					end
				end
			end
			else if (map[19:16] == 0 && map[23:20] > 0 && map[27:24] == 0 && map[31:28] == 0)
			begin
				map[31:28] <= map[23:20];
				if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
				begin
					map[23:20] <= 1;
				end
				else
				begin
					map[23:20] <= 0;
				end
			end
			else if (map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] == 0)
			begin
				map[31:28] <= map[27:24];
				map[27:24] <= 1;
			end
			else if (map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
			begin
			end
			else if (map[19:16] == 0 && map[23:20] > 0 && map[27:24] == 0 && map[31:28] > 0)
			begin
				if (map[31:28] == map[23:20])
				begin
					map[31:28] <= (map[31:28] + 1);
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
				else
				begin
					map[27:24] <= map[23:20];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
			end
			else if (map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0)
			begin
				if (map[27:24] == map[31:28])
				begin
					map[31:28] <= (map[31:28] + 1);
					map[27:24] <= 1;
				end
			end
			else if (map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] == 0)
			begin
				if (map[23:20] == map[27:24])
				begin
					map[31:28] <= (map[27:24] + 1);
					map[27:24] <= 0;
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
				else
				begin
					map[31:28] <= map[27:24];
					map[27:24] <= map[23:20];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
			end
			else if (map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0)
			begin
				if (map[31:28] == map[27:24])
				begin
					map[31:28] <= (map[27:24] + 1);
					map[27:24] <= map[23:20];
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
				else
				if (map[27:24] == map[23:20])
				begin
					map[27:24] <= (map[27:24] + 1);
					if ((map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0
				&& map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || (map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
				(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || (map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0))
					begin
						map[23:20] <= 1;
					end
					else
					begin
						map[23:20] <= 0;
					end
				end
			end
			else if (map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0)
			begin
			end

			/*Third line*/			
			
			if (map[35:32] > 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0)
			begin
				map[47:44] <= map[35:32];
				if 
				( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
				begin
					map[35:32] <= 1;
				end
				else
				begin
					map[35:32] <= 0;
				end
			end
			else if (map[35:32] > 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
			begin
				if (map[47:44] == map[35:32])
				begin
					map[47:44] <= (map[35:32] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
				else
				begin
					map[43:40] <= map[35:32];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
			end
			else if (map[35:32] > 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] == 0)
			begin
				if (map[43:40] == map[35:32])
				begin
					map[47:44] <= (map[35:32] + 1);
					map[35:32] <= 0;
					map[43:40] <= 1;
				end
				else
				begin
					map[47:44] <= map[43:40];
					map[43:40] <= map[35:32];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
			end
			else if (map[35:32] > 0 && map[39:36] > 0 && map[43:40] == 0 && map[47:44] == 0)
			begin
				if (map[39:36] == map[35:32])
				begin
					map[47:44] <= (map[35:32] + 1);
					map[35:32] <= 0;
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
					   	map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
				else
				begin
					map[47:44] <= map[39:36];
					map[43:40] <= map[35:32];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
					map[35:32] <= 0;
				end
			end
			else if (map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] == 0)
			begin
				if (map[43:40] == map[39:36])
				begin
					map[47:44] <= (map[43:40] + 1);
					map[43:40] <= map[35:32];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
					map[39:36] <= 0;
				end
				else
				if (map[35:32] == map[39:36])
				begin
					map[47:44] <= map[43:40];
					map[43:40] <= (map[39:36] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
					map[39:36] <= 0;
				end
				else
				begin
					map[47:44] <= map[43:40];
					map[43:40] <= map[39:36];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
					map[39:36] <= map[35:32];
				end
			end
			else if (map[35:32] > 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0)
			begin
				if (map[43:40] == map[47:44])
				begin
					map[47:44] <= (map[47:44] + 1);
					map[43:40] <= map[35:32];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
					    map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
					map[35:32] <= 0;
				end
				else
				if (map[35:32] == map[43:40])
				begin
					map[43:40] <= (map[43:40] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
				else
				begin
					map[39:36] <= map[35:32];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
			end
			else if (map[35:32] > 0 && map[39:36] > 0 && map[43:40] == 0 && map[47:44] > 0)
			begin
				if (map[39:36] == map[47:44])
				begin
					map[47:44] <= (map[47:44] + 1);
					map[43:40] <= map[35:32];
					map[39:36] <= 0;
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
				else
				if (map[35:32] == map[39:36])
				begin
					map[43:40] <= (map[39:36] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
					map[39:36] <= 0;
				end
				else
				begin
					map[43:40] <= map[39:36];
					map[39:36] <= map[35:32];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
			end
			else if (map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0)
			begin
				if (map[43:40] == map[47:44])
				begin
					map[47:44] <= (map[47:44] + 1);
					if (map[35:32] == map[39:36])
					begin
						map[43:40] <= (map[39:36] + 1);
						if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
						begin
							map[35:32] <= 1;
						end
						else
						begin
							map[35:32] <= 0;
						end
						map[39:36] <= 0;
					end
					else
					begin
						map[43:40] <= map[39:36];
						if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
						begin
							map[35:32] <= 1;
						end
						else
						begin
							map[35:32] <= 0;
						end
						map[39:36] <= map[35:32];
					end
				end
				else
				if (map[39:36] == map[43:40])
				begin
					map[43:40] <= (map[43:40] + 1);
					map[39:36] <= map[35:32];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
				else
				if (map[35:32] == map[39:36])
				begin
					map[39:36] <= (map[39:36] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[35:32] <= 1;
					end
					else
					begin
						map[35:32] <= 0;
					end
				end
			end
			else if (map[35:32] == 0 && map[39:36] > 0 && map[43:40] == 0 && map[47:44] == 0)
			begin
				map[47:44] <= map[39:36];
				if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
				begin
					map[39:36] <= 1;
				end
				else
				begin
					map[39:36] <= 0;
				end
			end
			else if (map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] == 0)
			begin
				map[47:44] <= map[43:40];
				map[43:40] <= 1;
			end
			else if (map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
			begin
			end
			else if (map[35:32] == 0 && map[39:36] > 0 && map[43:40] == 0 && map[47:44] > 0)
			begin
				if (map[47:44] == map[39:36])
				begin
					map[47:44] <= (map[47:44] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
				else
				begin
					map[43:40] <= map[39:36];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
			end
			else if (map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0)
			begin
				if (map[43:40] == map[47:44])
				begin
					map[47:44] <= (map[47:44] + 1);
					map[43:40] <= 1;
				end
			end
			else if (map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] == 0)
			begin
				if (map[39:36] == map[43:40])
				begin
					map[47:44] <= (map[43:40] + 1);
					map[43:40] <= 0;
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
				else
				begin
					map[47:44] <= map[43:40];
					map[43:40] <= map[39:36];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
			end
			else if (map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0)
			begin
				if (map[47:44] == map[43:40])
				begin
					map[47:44] <= (map[43:40] + 1);
					map[43:40] <= map[39:36];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
				else
				if (map[43:40] == map[39:36])
				begin
					map[43:40] <= (map[43:40] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
				)	
					begin
						map[39:36] <= 1;
					end
					else
					begin
						map[39:36] <= 0;
					end
				end
			end
			else if (map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0)
			begin
			end

			/*Forth line*/			
			
			if (map[51:48] > 0 && map[55:52] == 0 && map[59:56] == 0 && map[63:60] == 0)
			begin
				map[63:60] <= map[51:48];
				if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
				begin
					map[51:48] <= 1;
				end
				else
				begin
					map[51:48] <= 0;
				end
			end
			else if (map[51:48] > 0 && map[55:52] == 0 && map[59:56] == 0 && map[63:60] > 0)
			begin
				if (map[63:60] == map[51:48])
				begin
					map[63:60] <= (map[51:48] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
				else
				begin
					map[59:56] <= map[51:48];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] > 0 && map[55:52] == 0 && map[59:56] > 0 && map[63:60] == 0)
			begin
				if (map[59:56] == map[51:48])
				begin
					map[63:60] <= (map[51:48] + 1);
					map[51:48] <= 0;
					map[59:56] <= 1;
				end
				else
				begin
					map[63:60] <= map[59:56];
					map[59:56] <= map[51:48];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] > 0 && map[55:52] > 0 && map[59:56] == 0 && map[63:60] == 0)
			begin
				if (map[55:52] == map[51:48])
				begin
					map[63:60] <= (map[51:48] + 1);
					map[51:48] <= 0;
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
					   	map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
				else
				begin
					map[63:60] <= map[55:52];
					map[59:56] <= map[51:48];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
					map[51:48] <= 0;
				end
			end
			else if (map[51:48] > 0 && map[55:52] > 0 && map[59:56] > 0 && map[63:60] == 0)
			begin
				if (map[59:56] == map[55:52])
				begin
					map[63:60] <= (map[59:56] + 1);
					map[59:56] <= map[51:48];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
					map[55:52] <= 0;
				end
				else
				if (map[51:48] == map[55:52])
				begin
					map[63:60] <= map[59:56];
					map[59:56] <= (map[55:52] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
					map[55:52] <= 0;
				end
				else
				begin
					map[63:60] <= map[59:56];
					map[59:56] <= map[55:52];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
					map[55:52] <= map[51:48];
				end
			end
			else if (map[51:48] > 0 && map[55:52] == 0 && map[59:56] > 0 && map[63:60] > 0)
			begin
				if (map[59:56] == map[63:60])
				begin
					map[63:60] <= (map[63:60] + 1);
					map[59:56] <= map[51:48];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
					    map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
					map[51:48] <= 0;
				end
				else
				if (map[51:48] == map[59:56])
				begin
					map[59:56] <= (map[59:56] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
				else
				begin
					map[55:52] <= map[51:48];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] > 0 && map[55:52] > 0 && map[59:56] == 0 && map[63:60] > 0)
			begin
				if (map[55:52] == map[63:60])
				begin
					map[63:60] <= (map[63:60] + 1);
					map[59:56] <= map[51:48];
					map[55:52] <= 0;
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
				else
				if (map[51:48] == map[55:52])
				begin
					map[59:56] <= (map[55:52] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
					map[55:52] <= 0;
				end
				else
				begin
					map[59:56] <= map[55:52];
					map[55:52] <= map[51:48];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] > 0 && map[55:52] > 0 && map[59:56] > 0 && map[63:60] > 0)
			begin
				if (map[59:56] == map[63:60])
				begin
					map[63:60] <= (map[63:60] + 1);
					if (map[51:48] == map[55:52])
					begin
						map[59:56] <= (map[55:52] + 1);
						if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
						begin
							map[51:48] <= 1;
						end
						else
						begin
							map[51:48] <= 0;
						end
						map[55:52] <= 0;
					end
					else
					begin
						map[59:56] <= map[55:52];
						if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
						begin
							map[51:48] <= 1;
						end
						else
						begin
							map[51:48] <= 0;
						end
						map[55:52] <= map[51:48];
					end
				end
				else
				if (map[55:52] == map[59:56])
				begin
					map[59:56] <= (map[59:56] + 1);
					map[55:52] <= map[51:48];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
				else
				if (map[51:48] == map[55:52])
				begin
					map[55:52] <= (map[55:52] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[51:48] <= 1;
					end
					else
					begin
						map[51:48] <= 0;
					end
				end
			end
			else if (map[51:48] == 0 && map[55:52] > 0 && map[59:56] == 0 && map[63:60] == 0)
			begin
				map[63:60] <= map[55:52];
				if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
				begin
					map[55:52] <= 1;
				end
				else
				begin
					map[55:52] <= 0;
				end
			end
			else if (map[51:48] == 0 && map[55:52] == 0 && map[59:56] > 0 && map[63:60] == 0)
			begin
				map[63:60] <= map[59:56];
				map[59:56] <= 1;
			end
			else if (map[51:48] == 0 && map[55:52] == 0 && map[59:56] == 0 && map[63:60] > 0)
			begin
			end
			else if (map[51:48] == 0 && map[55:52] > 0 && map[59:56] == 0 && map[63:60] > 0)
			begin
				if (map[63:60] == map[55:52])
				begin
					map[63:60] <= (map[63:60] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
				else
				begin
					map[59:56] <= map[55:52];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
			end
			else if (map[51:48] == 0 && map[55:52] == 0 && map[59:56] > 0 && map[63:60] > 0)
			begin
				if (map[59:56] == map[63:60])
				begin
					map[63:60] <= (map[63:60] + 1);
					map[59:56] <= 1;
				end
			end
			else if (map[51:48] == 0 && map[55:52] > 0 && map[59:56] > 0 && map[63:60] == 0)
			begin
				if (map[55:52] == map[59:56])
				begin
					map[63:60] <= (map[59:56] + 1);
					map[59:56] <= 0;
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
				else
				begin
					map[63:60] <= map[59:56];
					map[59:56] <= map[55:52];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
			end
			else if (map[51:48] == 0 && map[55:52] > 0 && map[59:56] > 0 && map[63:60] > 0)
			begin
				if (map[63:60] == map[59:56])
				begin
					map[63:60] <= (map[59:56] + 1);
					map[59:56] <= map[55:52];
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
				else
				if (map[59:56] == map[55:52])
				begin
					map[59:56] <= (map[59:56] + 1);
					if ( 
					( 
						(map[3:0] > 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[3:0] != map[7:4] && map[7:4] != map[11:8] && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] == 0) || 
						(map[3:0] == 0 && map[7:4] > 0 && map[11:8] > 0 && map[15:12] > 0 && map[7:4] != map[11:8] && map[11:8] != map[15:12]) ||
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] > 0 && map[15:12] > 0 && map[11:8] != map[15:12]) || 
						(map[3:0] == 0 && map[7:4] == 0 && map[11:8] == 0 && map[15:12] > 0)
					)
					&& 
					(
						(map[19:16] > 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[19:16] != map[23:20] && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] == 0) || 
						(map[19:16] == 0 && map[23:20] > 0 && map[27:24] > 0 && map[31:28] > 0 && map[23:20] != map[27:24] && map[27:24] != map[31:28]) ||
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] > 0 && map[31:28] > 0 && map[27:24] != map[31:28]) || 
						(map[19:16] == 0 && map[23:20] == 0 && map[27:24] == 0 && map[31:28] > 0)
					)
					&& 
					(	
						(map[35:32] > 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[35:32] != map[39:36] && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] == 0) || 
						(map[35:32] == 0 && map[39:36] > 0 && map[43:40] > 0 && map[47:44] > 0 && map[39:36] != map[43:40] && map[43:40] != map[47:44]) ||
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] > 0 && map[47:44] > 0 && map[43:40] != map[47:44]) || 
						(map[35:32] == 0 && map[39:36] == 0 && map[43:40] == 0 && map[47:44] > 0)
					)
				)
					begin
						map[55:52] <= 1;
					end
					else
					begin
						map[55:52] <= 0;
					end
				end
			end
			else if (map[51:48] == 0 && map[55:52] == 0 && map[59:56] == 0 && map[63:60] == 0)
			begin
			end
		end
	end

endmodule
