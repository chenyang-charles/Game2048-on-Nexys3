`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    22:35:29 01/04/2015 
// Design Name: 
// Module Name:    number 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module number(
			input wire clka,
			input wire [15:0] addra,
			output reg douta
    );

	parameter data = {
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000011111111100000000000000000000000000000,
70'b0000000000000000000000000000111111111111111000000000000000000000000000,
70'b0000000000000000000000000011111111111111111100000000000000000000000000,
70'b0000000000000000000000001111111111111111111110000000000000000000000000,
70'b0000000000000000000000011111111111000011111110000000000000000000000000,
70'b0000000000000000000000111111111000000000111110000000000000000000000000,
70'b0000000000000000000000111111000000000000011110000000000000000000000000,
70'b0000000000000000000000111100000000000000011110000000000000000000000000,
70'b0000000000000000000000010000000000000000111110000000000000000000000000,
70'b0000000000000000000000000000000000000000111110000000000000000000000000,
70'b0000000000000000000000000000000000000001111100000000000000000000000000,
70'b0000000000000000000000000000000000000011111100000000000000000000000000,
70'b0000000000000000000000000000000000000011111000000000000000000000000000,
70'b0000000000000000000000000000000000000111111000000000000000000000000000,
70'b0000000000000000000000000000000000001111110000000000000000000000000000,
70'b0000000000000000000000000000000000001111100000000000000000000000000000,
70'b0000000000000000000000000000000000011111100000000000000000000000000000,
70'b0000000000000000000000000000000000111111000000000000000000000000000000,
70'b0000000000000000000000000000000001111110000000000000000000000000000000,
70'b0000000000000000000000000000000011111100000000000000000000000000000000,
70'b0000000000000000000000000000000011111100000000000000000000000000000000,
70'b0000000000000000000000000000000111111000000000000000000000000000000000,
70'b0000000000000000000000000000001111110000000000000000000000000000000000,
70'b0000000000000000000000000000011111100000000000000000000000000000000000,
70'b0000000000000000000000000000011111000000000000000000000000000000000000,
70'b0000000000000000000000000000111111000000000000000000000000000000000000,
70'b0000000000000000000000000001111110000000000000000000000000000000000000,
70'b0000000000000000000000000001111111111111111100000000000000000000000000,
70'b0000000000000000000000000011111111111111111100000000000000000000000000,
70'b0000000000000000000000000011111111111111111100000000000000000000000000,
70'b0000000000000000000000000001111111111111111100000000000000000000000000,
70'b0000000000000000000000000000000000111110000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000011110000000000000000000000000000000000000,
70'b0000000000000000000000000000011111000000000000000000000000000000000000,
70'b0000000000000000000000000000111110000000000000000000000000000000000000,
70'b0000000000000000000000000000111110000000000000000000000000000000000000,
70'b0000000000000000000000000001111100000000000000000000000000000000000000,
70'b0000000000000000000000000001111100000000000000000000000000000000000000,
70'b0000000000000000000000000011111000000000000000000000000000000000000000,
70'b0000000000000000000000000011111000000011110000000000000000000000000000,
70'b0000000000000000000000000011111000000011110000000000000000000000000000,
70'b0000000000000000000000000111110000000011110000000000000000000000000000,
70'b0000000000000000000000000111110000000011110000000000000000000000000000,
70'b0000000000000000000000001111100000000011110000000000000000000000000000,
70'b0000000000000000000000001111100000000011110000000000000000000000000000,
70'b0000000000000000000000001111100000000011110000000000000000000000000000,
70'b0000000000000000000000011111000000000111110000000000000000000000000000,
70'b0000000000000000000000011111000000000111110000000000000000000000000000,
70'b0000000000000000000000011111000000000111110000000000000000000000000000,
70'b0000000000000000000000111110000000000111110000000000000000000000000000,
70'b0000000000000000000000111110000000000111110000000000000000000000000000,
70'b0000000000000000000000111110000000000111110000000000000000000000000000,
70'b0000000000000000000000111110000000000111110000000000000000000000000000,
70'b0000000000000000000000111111111111111111111111110000000000000000000000,
70'b0000000000000000000000111111111111111111111111110000000000000000000000,
70'b0000000000000000000000111111111111111111111111110000000000000000000000,
70'b0000000000000000000000111111111111111111111111100000000000000000000000,
70'b0000000000000000000000000011111111111111110000000000000000000000000000,
70'b0000000000000000000000000000000000000011110000000000000000000000000000,
70'b0000000000000000000000000000000000000011110000000000000000000000000000,
70'b0000000000000000000000000000000000000011110000000000000000000000000000,
70'b0000000000000000000000000000000000000011110000000000000000000000000000,
70'b0000000000000000000000000000000000000011110000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000111100000000000000000000000000000000,
70'b0000000000000000000000000000011111111111110000000000000000000000000000,
70'b0000000000000000000000000001111111111111111100000000000000000000000000,
70'b0000000000000000000000000011111111111111111111000000000000000000000000,
70'b0000000000000000000000000011111111101111111111000000000000000000000000,
70'b0000000000000000000000000111111000000000111111000000000000000000000000,
70'b0000000000000000000000000111110000000000001110000000000000000000000000,
70'b0000000000000000000000000111100000000000000000000000000000000000000000,
70'b0000000000000000000000000111100000000000000000000000000000000000000000,
70'b0000000000000000000000000111100000000000000011000000000000000000000000,
70'b0000000000000000000000000111110000000000011111000000000000000000000000,
70'b0000000000000000000000000111111000000011111111100000000000000000000000,
70'b0000000000000000000000000111111100001111111111100000000000000000000000,
70'b0000000000000000000000000011111110111111111110000000000000000000000000,
70'b0000000000000000000000000001111111111111110000000000000000000000000000,
70'b0000000000000000000000000000111111111111000000000000000000000000000000,
70'b0000000000000000000000000000011111111110000000000000000000000000000000,
70'b0000000000000000000000000000111111111111100000000000000000000000000000,
70'b0000000000000000000000000001111111111111110000000000000000000000000000,
70'b0000000000000000000000000011111110011111111000000000000000000000000000,
70'b0000000000000000000000000011111100000111111100000000000000000000000000,
70'b0000000000000000000000000111111000000011111100000000000000000000000000,
70'b0000000000000000000000000111110000000000111110000000000000000000000000,
70'b0000000000000000000000000111110000000000111110000000000000000000000000,
70'b0000000000000000000000000111100000000000011110000000000000000000000000,
70'b0000000000000000000000000111100000000000111110000000000000000000000000,
70'b0000000000000000000000000111110000000000111110000000000000000000000000,
70'b0000000000000000000000000111111000000001111110000000000000000000000000,
70'b0000000000000000000000000011111111000111111100000000000000000000000000,
70'b0000000000000000000000000011111111111111111100000000000000000000000000,
70'b0000000000000000000000000000111111111111111000000000000000000000000000,
70'b0000000000000000000000000000011111111111100000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000011111100000000000000,
70'b0000000000000000000000000000000000000000000000011111111111100000000000,
70'b0000000000000000000000000000000000000000000001111111111111000000000000,
70'b0000000000000000000000000000000000000000000111110001111110000000000000,
70'b0000000000000000000000000000000000000000001111000000001100000000000000,
70'b0000000000000000000000000000000000000000011100000000000000000000000000,
70'b0000000000000000000000001100000000000000111000000000000000000000000000,
70'b0000000000000000000000011100000000000001111000000000000000000000000000,
70'b0000000000000000000001111100000000000011110000000000000000000000000000,
70'b0000000000000000000111111100000000000011100000000000000000000000000000,
70'b0000000000000000011111111100000000000111100000000000000000000000000000,
70'b0000000000000001111111111000000000001111100000000000000000000000000000,
70'b0000000000000001111001111000000000001111000000000000000000000000000000,
70'b0000000000000001110001111000000000001111000011111111000000000000000000,
70'b0000000000000000000001111000000000011111001111111111100000000000000000,
70'b0000000000000000000001111000000000011110011111111111110000000000000000,
70'b0000000000000000000001111000000000011110111100011111110000000000000000,
70'b0000000000000000000001111000000000011111110000000111111000000000000000,
70'b0000000000000000000011111000000000111111100000000011111000000000000000,
70'b0000000000000000000011111000000000111111000000000011111000000000000000,
70'b0000000000000000000011110000000000111111000000000001111000000000000000,
70'b0000000000000000000011110000000000111110000000000001111000000000000000,
70'b0000000000000000000011110000000000111110000000000001111000000000000000,
70'b0000000000000000000011110000000000011111000000000001110000000000000000,
70'b0000000000000000000011110000000000011111000000000001110000000000000000,
70'b0000000000000000000011110000000000011111100000000011100000000000000000,
70'b0000000000000000000011110000000000001111100000000111100000000000000000,
70'b0000000000000000000111110000000000001111111000001111000000000000000000,
70'b0000000000000001111111111111100000000111111111111110000000000000000000,
70'b0000000000000111111111111111000000000011111111111100000000000000000000,
70'b0000000000000111111111111110000000000001111111110000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000111110000000000000000001111100000000000000000000,
70'b0000000000000000000111111111100000000000001111111111000000000000000000,
70'b0000000000000000011111111111110000000001111111111111110000000000000000,
70'b0000000000000000111100001111111000000011111111111111110000000000000000,
70'b0000000000000000110000000111111000000111100000011111111000000000000000,
70'b0000000000000000000000000011111000000110000000000111111000000000000000,
70'b0000000000000000000000000011111000000000000000000111111000000000000000,
70'b0000000000000000000000000011111000000000000000000011111000000000000000,
70'b0000000000000000000000000011110000000000000000000011111000000000000000,
70'b0000000000000000000000000111110000000000000000000011111000000000000000,
70'b0000000000000000000000000111100000000000000000000011110000000000000000,
70'b0000000000000000000000011111000000000000000000000011110000000000000000,
70'b0000000000000000000001111100000000000000000000000111100000000000000000,
70'b0000000000000000011111110000000000000000000000001111000000000000000000,
70'b0000000000000000111111111110000000000000000000001110000000000000000000,
70'b0000000000000001111111111111000000000000000000011100000000000000000000,
70'b0000000000000001111111111111100000000000000000111000000000000000000000,
70'b0000000000000000000000111111110000000000000011110000000000000000000000,
70'b0000000000000000000000001111110000000000000111100000000000000000000000,
70'b0000000000000000000000000111110000000000111111000000000000000000000000,
70'b0000000000000000000000000011110000000111111100000000000000000000000000,
70'b0000000000000000000000000011110000001111111111111111111000000000000000,
70'b0000000000000000000000000011110000011111111111111111111000000000000000,
70'b0000000000000000000000000011110000111111111111111111110000000000000000,
70'b0000000000000000000000000011100000000011111111111111100000000000000000,
70'b0000000000000000000000000111100000000000000000000000000000000000000000,
70'b0000000000000000000000001111000000000000000000000000000000000000000000,
70'b0000000000000111100000011110000000000000000000000000000000000000000000,
70'b0000000000001111111111111100000000000000000000000000000000000000000000,
70'b0000000000011111111111110000000000000000000000000000000000000000000000,
70'b0000000000011111111111000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000001111110000000000000000000000000000000000000,
70'b0000000000000000000000001111111111110000000000000000000000000000000000,
70'b0000000000000000000000111111111111100000000000000000000000000000000000,
70'b0000000000000000000011111100111111000000000000000000000000000000000000,
70'b0000000000000000000111100000000110000000000000000000000000000000000000,
70'b0000000000000000001110000000000000000000000000000000000000000000000000,
70'b0000000000000000011100000000000000000000000000000000000010000000000000,
70'b0000000000000000111100000000000000000000000000000000000110000000000000,
70'b0000000000000001111000000000000000000000000000000000001110000000000000,
70'b0000000000000011110000000000000000000000000000000000111110000000000000,
70'b0000000000000011110000000000000000000000000000000001111110000000000000,
70'b0000000000000111100000000000000000000000000000000011111110000000000000,
70'b0000000000000111100000000000000000000000000000000111111110000000000000,
70'b0000000000001111100001111111100000000000000000001111111110000000000000,
70'b0000000000001111000111111111110000000000000000011111111110000000000000,
70'b0000000000001111001111111111111000000000000000111110111100000000000000,
70'b0000000000001111011110001111111000000000000001111100111100000000000000,
70'b0000000000011111111000000111111000000000000011110000111100000000000000,
70'b0000000000011111110000000011111100000000000111100000111100000000000000,
70'b0000000000011111100000000001111100000000001111000000111100000000000000,
70'b0000000000011111100000000001111100000000011110000000111100000000000000,
70'b0000000000011111000000000000111100000000111100000001111100000000000000,
70'b0000000000011111000000000000111000000001111000000001111100000000000000,
70'b0000000000011111100000000000111000000011110000000001111100000000000000,
70'b0000000000001111100000000001111000000111111100000001111000000000000000,
70'b0000000000001111100000000001110000001111111111111111111000000000000000,
70'b0000000000001111110000000011110000111111111111111111111111111000000000,
70'b0000000000000111111000000111100000111111111111111111111111110000000000,
70'b0000000000000011111111111111000000000000000111111111111111100000000000,
70'b0000000000000001111111111110000000000000000000000001111111000000000000,
70'b0000000000000000111111111000000000000000000000000001111000000000000000,
70'b0000000000000000000000000000000000000000000000000011111000000000000000,
70'b0000000000000000000000000000000000000000000000000011111000000000000000,
70'b0000000000000000000000000000000000000000000000000011110000000000000000,
70'b0000000000000000000000000000000000000000000000000011110000000000000000,
70'b0000000000000000000000000000000000000000000000000011110000000000000000,
70'b0000000000000000000000000000000000000000000000000011110000000000000000,
70'b0000000000000000000000000000000000000000000000000010000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000111111100000000000,
70'b0000000000000000000000000000000000000000000000000011111111110000000000,
70'b0000000000000000000000000000000000000000000000000111000111110000000000,
70'b0000000000000000000000000000000000000000000000001110000011111000000000,
70'b0000000000000000000100000000000000000000000000001110000001111000000000,
70'b0000000000000000011100000000000111111110000000001110000001111000000000,
70'b0000000000000001111100000000011111111111000000001111000001110000000000,
70'b0000000000000111111100000000111111111111100000001111100001110000000000,
70'b0000000000011111111100000001110000011111100000001111110011100000000000,
70'b0000000000011110111000000000000000001111100000000111111111000000000000,
70'b0000000000011000111000000000000000000111100000000011111110000000000000,
70'b0000000000000000111000000000000000000111100000000111111110000000000000,
70'b0000000000000000111000000000000000000111100000001111111111100000000000,
70'b0000000000000001111000000000000000000111000000011110001111100000000000,
70'b0000000000000001111000000000000000001111000000111100000111110000000000,
70'b0000000000000001111000000000000000001110000000111000000011110000000000,
70'b0000000000000001111000000000000000011100000001111000000011110000000000,
70'b0000000000000001111000000000000001111000000001111000000001110000000000,
70'b0000000000000001110000000000000011110000000001111000000001110000000000,
70'b0000000000000001110000000000001111100000000001111100000011110000000000,
70'b0000000000000001110000000001111110000000000001111110000011100000000000,
70'b0000000000011111111111000011111111111111100000111111111111000000000000,
70'b0000000000111111111111000111111111111111100000011111111110000000000000,
70'b0000000000111111111110000111111111111111000000001111111000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000001111111000000,
70'b0000000000000000000000000000000000000000000000000000000111111111100000,
70'b0000000000000000000000000000000000000000000000000000011111111111000000,
70'b0000000000000000000000000000000000000000000000000000111000000110000000,
70'b0000000000000000000000000000000000000000000000000001110000000000000000,
70'b0000000000000001111110000000000000000000000000000011100000000000000000,
70'b0000000000001111111111100000000011111111111100000111000000000000000000,
70'b0000000000011111111111100000000111111111111000001111000000000000000000,
70'b0000000000111000001111110000001111111111110000001110000000000000000000,
70'b0000000000110000000111110000001110000000000000011110000000000000000000,
70'b0000000000000000000011110000001110000000000000011110011111110000000000,
70'b0000000000000000000011110000001110000000000000011100111111111000000000,
70'b0000000000000000000011110000001110000000000000111111111111111100000000,
70'b0000000000000000000011100000011110000000000000111111000001111100000000,
70'b0000000000000000000111100000011111111000000000111110000000111100000000,
70'b0000000000000000001111000000011111111110000000111110000000111100000000,
70'b0000000000000000001110000000011111111111000000111100000000011100000000,
70'b0000000000000000011100000000000000111111100000111100000000011100000000,
70'b0000000000000001111000000000000000001111100000111110000000011100000000,
70'b0000000000000111110000000000000000000111100000111110000000111000000000,
70'b0000000000011111000000000000000000000011100000011111000000111000000000,
70'b0000000001111111111111110000000000000011100000011111100011110000000000,
70'b0000000011111111111111110000000000000011100000001111111111100000000000,
70'b0000000111111111111111100000000000000011100000000111111110000000000000,
70'b0000000000000000000000000000000000000111000000000000000000000000000000,
70'b0000000000000000000000000000000000001111000000000000000000000000000000,
70'b0000000000000000000000000000111110111110000000000000000000000000000000,
70'b0000000000000000000000000001111111111000000000000000000000000000000000,
70'b0000000000000000000000000011111111110000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000001100000000000000000000000000000000,
70'b0000000000000000001111111111000000011100000000011111111000000000000000,
70'b0000000000000000011111111110000000111100000000111111111100000000000000,
70'b0000000000000000111111111110000011111100000001111011111110000000000000,
70'b0000000000000000111000000000001111111100000001100000111110000000000000,
70'b0000000000000000111000000000001110111100000000000000011110000000000000,
70'b0000000000000000111000000000001100111100000000000000011110000000000000,
70'b0000000000000001110000000000000000111000000000000000011110000000000000,
70'b0000000000000001110000000000000000111000000000000000011110000000000000,
70'b0000000000000001111110000000000000111000000000000000011100000000000000,
70'b0000000000000001111111100000000000111000000000000000111000000000000000,
70'b0000000000000001111111110000000000111000000000000000111000000000000000,
70'b0000000000000001111111111000000000111000000000000001110000000000000000,
70'b0000000000000000000011111000000000111000000000000011100000000000000000,
70'b0000000000000000000000111100000001111000000000001111000000000000000000,
70'b0000000000000000000000111100000001111000000000011110000000000000000000,
70'b0000000000000000000000011100000001111000000011111100000000000000000000,
70'b0000000000000000000000011100001111111111000111111111111110000000000000,
70'b0000000000000000000000011000011111111111001111111111111110000000000000,
70'b0000000000000000000000011000011111111110001111111111111100000000000000,
70'b0000000000000000000000111000000000000000000000000000000000000000000000,
70'b0000000000000011000001110000000000000000000000000000000000000000000000,
70'b0000000000000111111111100000000000000000000000000000000000000000000000,
70'b0000000000001111111111000000000000000000000000000000000000000000000000,
70'b0000000000000111111100000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000001000000000000000000000000000011000000000000000000000000110000,
70'b0000000111000000000000011111100000000011111100000000000000000001110000,
70'b0000001111000000000001111111111000000011111110000000000000000011110000,
70'b0000011111000000000111111111111100000001111111000000000000000011110000,
70'b0000111111000000001111110001111110000000001111100000000000000111110000,
70'b0001111111000000001111000000011110000000000111110000000000001111110000,
70'b0011111111000000011110000000001111000000000011110000000000011111110000,
70'b0011110111000000011110000000001111000000000001110000000000011111110000,
70'b0001100111000000011100000000000111000000000001110000000000111111110000,
70'b0000000111000000011100000000000111000000000011110000000001111011110000,
70'b0000000111000000011100000000000111000000000011110000000011110011110000,
70'b0000000111000000011100000000001111000000000111100000000111100011110000,
70'b0000000111000000011110000000001111000000001111100000000111100011110000,
70'b0000000111000000011110000000001110000000001111000000001111111111111100,
70'b0000001111000000001111000000011110000000011110000000011111111111111100,
70'b0000001111000000001111100001111100000001111100000000000000000011110000,
70'b0000001111000000000111111111111100000011111000000000000000000011110000,
70'b0000001111000000000011111111111000000111111111111000000000000011110000,
70'b0000001111000000000000111111100000001111111111111000000000000011110000,
70'b0000000000000000000000000000000000001111111111111000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0001111000000000000000000000000000000000000000011000000000001111110000,
70'b0001111110000000000000011111110000000000000000111000000000111111111000,
70'b0001111111100000000000111111111100000000000000111000000001111111111100,
70'b0000011111110000000011111111111110000000000001111000000001111000111100,
70'b0000000011111000000011111000011111000000000011111000000001110000011110,
70'b0000000001111000000111100000001111100000000111111000000001110000011110,
70'b0000000000111000000111100000000111100000001111111000000001110000011110,
70'b0000000000111100001111000000000011100000001111111000000001111000111100,
70'b0000000000111100001111000000000011100000011110111000000001111111111100,
70'b0000000000111000001110000000000011100000111100111000000000111111111000,
70'b0000000001111000001110000000000011100001111000111000000000111111111100,
70'b0000000011111000001111000000000011100001111000111000000001111000111100,
70'b0000000011110000001111000000000111100011111111111111000001110000011110,
70'b0000000111100000000111100000000111100111111111111111000011110000011110,
70'b0000001111000000000111110000001111000111111111111111000011110000011110,
70'b0000011110000000000011111000111111000000000000111000000011110000011110,
70'b0001111101111110000011111111111110000000000000111000000001111000111100,
70'b0011111111111110000000111111111100000000000000111000000001111111111100,
70'b0111111111111110000000001111100000000000000000111000000000111111111000,
70'b0000000000000010000000000000000000000000000000000000000000001111100000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000,
70'b0000000000000000000000000000000000000000000000000000000000000000000000
};

	always @(posedge clka)
	begin
		douta <= data[53899 - addra];
	end

endmodule
